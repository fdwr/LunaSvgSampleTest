��  �bnnnnaWnnnnnnnnabbbabv�����vnaLOOOOWWWOLOLLOWOTavp�vnaOLLOW���ynnnv�����������������������vngaYaaavvnaanvz�yaaanaYOE4)%))=EEOOanbgp������v���������nappzz���vpaanvwnnpv��w��������wy�z���ppwpnv�����������n^aanaWEEEE=ELOOA46699OY\an���������ynWnnapvv�y�����������ż���������pbOajnbaWnaannnnnnv����yp���nbWbannnnnWbbnnnanvvvnW]]OOWbbn�������naOOE<DEO]OOOTWnnabnpp�vnaOD<DWv������v�����������������������vnvnaa]Wnvnnanp���waaWWOOO<,)%%)6=<EEOWbpy�����������������vrpv����zpagpzzvgapp�vpz�������wpvw���zvzv�������������nnwpaOLAAE666<A6)4669L^YYv����������vnnnpvp���������������Ũ�������pWWa]bWabnnnnnnnnnv���������nnbaannnnnOObnnnavyvaW]TOOOWan��������vnWDE<69<LW]]TTbnnnnppv�vnaEBBDOv���������������������������������n�nnnWnnnanyy���waYOWOEE6)#/7=<<EWbvz�����������������yzvpz�y�wpagn���nabgnpwz�������zvvv����z��������������������nWEAE6/,-//,%)446EOT\v������¨���vv�vvpv����������������Ϸ�������pWOOT]Waannnnnnanavy���������nnnannnnan<DbabnnvynaOWTOOObn�������yvnO<<<4.4<Wa]]WappyvvvnvnnaE<<DWv������������������ż��������������v�pnnnanaany����wWOOOEE?6%/=8<6ERbvz�������������������vpzzyzpvppn���paWWgnwz��������vvv��������������ż��������nRE<<4))-,%)69BLOav������ڱ������zvv�����������������˼��ż��ynOOObWWannnabbWb]nvyy�������nnnnnnnabb,<TWbnnvvnWOTOWWWbpy�������vnbO<<4/4/<OWTW]anvyyvvnnabWE99BOv�������������������ű������������v�nnnnnnnanz����waYOEE?E6/<6<6<Wnz���������������������y���pyvyv���vaYYagnvv�����zvvpw��������������ȼ¼������pWEB<-%%,%)/BTYn��������¤�������vv��������������������ų���nOETjWabnanabWWWannvy��������nnnnnnaaaa-EWb]WnvvaaOLW]aYnny�������vbO<</-,444ALWannpnyyvnabbaWOE<<Da�������������������¼����������vvvypnpnapwz������vaRHEOH6)+6EE=<HYv��������������������������wry�����pn^Y\a\gy�zzpvpg\mv����������������ż������aRE=/%,,%%-6Bnnv��������ѳ��������������������������ż�����nWOO]babbaabnWOT]]]nvy�������vnnnnnnnnan%9ELOWbnnaOLOabjjnny�������vWD<6/,,4/49DWanpyy�yyaOLOWWWOEDOWn��������������������˼��������vv����vv���������vaWEERY>))*)6DRPOEOav������������������������z�prw�������rnaOPSYapnpppnpnggh��������������������¨���pbH</%,%%-/<Onn�����������¼���v�������������������ż�����vnWT]anbWbWWWODLTTWbnv��vvvnnnnnnnnn/49DOannWDIIbnnnpp�������nbE<964.//9BWannv����nbLBOWaaWOWWbn�������������������ϳ��������vnv������wz��������paOEDHRE//6<EOaaaWOaw������������������������zrvwr�������waYE?EYgg\agg\aagrpy�������������������³��znnR</)46Oav�������������±������������������������ż�����aWLWnaaOOEE<9<DLOannn��vvvnnnnnnnnnnn6<E]nbOEBL]nvyy���nnnTD6<<<6/9EWannvy���vaTDOObnabWnnvv������������������ϼ����������zvn�����zzv�������wpWE>>DO=6<EER\pgnaWav�����������������z�����zwmzwz�������zaYE<??YWWYYaY\amrv��������������������ų��vpgR<,,6EWn���������������ϱ��������������������������ż�����vjTWabaOOOD946DLLOWWanvyvnnnnnnvnnaann%4<LWWOOOLWv����yvnaWTL<6),/46<DWnnnnvvyvvnbWWWbannnv�����������v���������ż���������nv����zvz����zypa[O</66<=DE?EWgzzwn\nv���yzz�����������w�����prnvv��������znYO???EOOYaYagarzz����������������¼������na[H</*<Eap���������������ڼ�������������������¹�����Ź�����naaWWOIBBD<4BEELDIDOWnnnnabbannnabbnn%.<LIDOWYbv����ypnbbOD<9/)%6<L]nnvvnnbWanaabnnvnnn���������������y��������������������yvvvzzz��v���pwnnaWO<6666/8??EOWv��ywnvpaaangr�����������������waggw���������rnYYYEEEOYaaapzz�������������������������wpgOD<))%)<Ony����������������ϼ����������������¹������¼�������ynWODD<BBBB<DLE<<96DWWWWWWabnnbbWWWW/4B<O]Ynv��nnaWOE94/))6DWnnypnpnWO]bnabvvvv������������vvz����������������������yrnnnnww���vkabWEE<6/+////<EOOYnvv�wpgaPOOYWam�����������������a\\n����������wmnYOOOannmrr����������zzv������������wggaR>6.#)9Wpz����������������ű�������������ϼ�����������¹�����nWI<B<DBIOOOLLB9449DLBDOWannbWWWWWO-6BEWnnv��pbanWOB4.6)./6Onvyvvypn]T]Tanv���������������yvv������������������������znannn���vaWOODD<6/*))%//=EOYagnpwraYPEE???Okw���������������wgYgzz����������wp\Y\nwwwrrw���������znan������������ygaaWRE6+*,=Oa���������������Ź�������������������������������������naD<6<DLT]]a]DEA94/99<BEOWanabWbWaa)4DOn������nnabWE<//6,%.9DWbvvyy�ynjbaabn����������ż�������v��������������������������znnvnpzzpgRE6666/)*<=<OYaargaa>666+/6Ean���������������p\Yhzrr���zz�����wrrz����zzz���������zmgw�����������vpY\RRRH<.),<Oaw����������������������������������������������������znWL666DOT]a]]WOE</,/6<DOOOWannanbbW
%-.<Wn������vnnbWOB644/),.<Waan����vnnvnv������������ϼ�������������������������������������wnnagO>9/+*)*)#26<EOYWWYWO=///+*/=OYp��z���������vn\a\mzrrwwzwz�������������������������zzz������������v[SORWROD6*/<WYpw�����yv�������������������������������������������vnWOA69EO]]nnnaj]B64.6<DEWWbnnnnnbbO
%)/6<Wv������vvaWOE96/-/,,4IOaanv�����vvn��������������ϼ��������������������vnvy�����������zaROE6./66=EEE<<<<//*/6<Raannpppz����rgY\ngmanngpr�������������������������������������z���aR?ERRRWE<6)%)+.<OWW]vvwvnnnnnv��������������������������������������ynWAE<OTbbnnnpnaWIB996BDOWbannnnnaWO
,-/./9av���vnnWOD63/,,).<DOany������vnn��������������Ź����������������vvvnnny�����������v[O?6/


)-//76/)*+$**/6?OOYYWaaprpwraY\\nnc\\Yaaaw�����������������������������������wwz�znYE=?WROEE<6/+#).6<DOOOWaa\WTLOOaaannvn������������������������������������pTDBLWbnvvvynWW]EE<ADOWannnnnaaWW,/,))6Wn��vvnvnnWOD66/,//<DDWavvyy���ynv����������������ϼ���������������nnnnaanzz���������p[RD6*
/.)*/6=EEEEWRgwaYWYWYYa\SRYWYaw�����������Ƽ������ż��������������zgagaYWE?OYWE?EE<D<4/..6<DE?<<?OOHLA=EEEOOEanv��������������������������yvbv��n]E<OWnpv����vbnaaWE<DObnnnnnabbWW
%4.)/On��nnnnnnnnWI<<63<DDWbnnvvpnvvvyyv�����������������®�������������nnnYWWYnn����������pWH<%#**7626<OO\nYE=POY\a\YHOYanz��������������������Ƽ�������������vaYROOSO?OYYOEOEEOO<6666<<6<6+.<DDE666===<BLWn������ż����������������zban�vvjTEObnnv����yvppnbTOOOanvvnnnnnWW
%6/-/Lnvyynnb]nnnbWEDBB<DWWbnvvnnanvnpy��v����������������³������Ź����vnnkaWWWnz�����������bG6))%$*/2/55EOW\PE==EWaaa\OO\avz������ƽƽ���������Ƽ��������������gaRE6HHOEOOOWSYROOWOE<<D6.#))).66696==6///=LTany�����������n���������vvznanbaannnnjYWWannp�������pnanbbbbnnnvnnnbn

,.6)4Obnyyvnn]]a]OTBDIBOOWWnvnpvnnvv��������������������ż�������¨���vnnnnaaYaanw�����������nD/
)	
)***//+225??EE=66=ParraPS\anw������ƽƽ���������ż�������������zg\R<6=EHEEE?ORa\WWWYWRRD6)#)).636A<644-/6=LTav����������v��������yvnWWbaWbannnnnananpy���v���ynnnnabbbbnnnnnnn%),))/LO]nppjbb]TL99<BLLIOObnv�vpvvvv������������������������¼��¼�����vvnaaannpnnnn������������a=)

*+/!!$!/**/26866===6=O\nmaY\gnvz���ý�����������ƽƽ��������������w\YO<56<=EE=EHR\pnWWOObWH</))).6=///4/66AAOkn�������ynvv�������pbnWWaWOWWnnpvynnpy�vy�nnnanabOOWWWWbbb.//,)9BOWbWWW]OD<4449DBLE]Wanvz��������������������������������·�����nnnYWYanvvvw�������������W=+%).//**!#&!//2$!**265=656=EEHOPYaaagzwz������������������ƽ�������������rwwp\R?<5/=?OEEEHEOavgWWOWWWO</).36///66AAOTWa^Wanv�����pnbv��������vvnbnbbaWWnv����vnpyvypnnnnvnnaa]]]TBDDOOOWbBD<6,%))/9<<IOWOOOLBB4,/46<ALTWabpy���vv��������������������������ŷ������pnYWOU^n����������������vWO76///)))%)66/2*!	)$!$/5=52/*/65E==6==HPaYYPYYgw�������������ƽ�����ƽ�������������wgmnnWR<82+<?OOEEEEOapp\O<OWWW=6).66//.6=BOWa^T<EOWnnnvngnabv�����������n]bbaWbanv�����vpynnaWOWnnnnnnYWLL9/6<DDOOnOOWB./4/66669DBDIDOLB<64/449LTa]bap�������������������������������Ѽ������n^LLLLar������������z��ppaO<=EEE6/#)%/6<7///!	**//6=EP?====?PPE==ERammaSYaz��������������ƽ�������������������zaY\naYOE5/*6=OP=?OOWannYYE=OWYO6+.)36<<<?EOYaTL<AOEPOOY\WWaan��������zypWTWWbbanz����znppnaWOELOananaYO<9.,46BObnWWOD99B<<<,-,9B9B<IOO<6649<BW]nnap�������������ŷ��������������������Ѽ�����nOE=AOav�����������v�vwggYE=EYWEO?6/)//6=?=6//	//226=EEPOHH?JPYaSEEHSahanYan�������������̼�������������zzz�����a\YYWOROP8//6=OO=EY\grmaYOEEOOOO?66/)).3<OEEEHEOOTA6AE=5=AEAEOWWWnnvv�vppnnWTOWWan����v]bjaOE9<EOObbnbWL9.),6DWbnnaOLTTWO</)-.9<<ADLO<<<BBTbjnvnp���������������ų��������������������Ź��aOA=ATnw�����������vnvpgYOE=WaaaWOE<<?<EHE<52**$/668?EHPYacYY\\hYYSOSYY\ahnmz����ƹ�������Ƽ����������zhmmggpz��z[SE=E<EEO=627EEEEPgnnnaRE?EYYWWOHOE<6)))#/<>OOOOOEEOYOBEE=6///-6=EOOOWbnvnnvvvnaWbTOWav����aW]aWL<4<OLT]abbOA-),4EOWvnbW]nnWD9,)46ELOTWOEBEEWanpnv������������������¨������������������Ἠ��vaYEEETnz����������vggnbYWWEHYrwrpaa\\YYOEE62*+*/!+5==EHHEOYhraga\\SYaYY\\S\aar�����ý������������������waYY\\\agnp\FEE===?JOO==<EEHRWgnnnaP?HSYanaWWWWWH6/..<>HHDOOOOEOWOOE<//)%)/9DOIIOOaanvvvvbW]TWIWbnz���vaTTTOB<9BDTT]aaE<<,))69LW�ynabnnbW<4-/9ETYaTLOWWWWapvvv�������������������ų������������������Ϲ����pnaOUYknw����������vnggYRYaYYgz���wwrwnnOE7//#*//*!/?=??HOOYSagrmnaY\Yc\YYa\\\\cr�����ýƳ�������������zwmcYYSYYa\ccSJEEEE=5EEOYROPE??Ra\gWaY\OOPanaaanaaYWE<<<>DD>RWWOOEOYaYO</%-4B<<<IOWannvvnnWWWabnnnnz�nOTWD9BBLOTTbaW<96/49BTWvynnnnvnW</,,6BWaaWOYnnnnnv���������������������¼�����������������ڼ�����yvvavwpw����������vvvaSS\nrmzz���z���vaR<6//65562**//=PPYORY\hnmw�wmaYY\aaarng\\\hnz�������������������wzrwaYOYPSahaSOHEEOEE?58?OYgaYEEORaaaEORaY\Ya^gapnpgnbWOGHODHOOOOEOOSWYaLA/--//.6<DOOWnvnnvnnvaannapyynaWOLA9<LTOTTTTOO6,)-6BLWWnnyvyvvvnO<66469EWWWWnvvnv�����������������������¼�ż��������������ų�����������vpzy���������yvvYYYp���zwzzw��zngS=///6==?825?=OOYYgahgwrrrwrwraYYahmmrhh\aacrz�������������zwwwwwwzwmmaYOPS\aYRE=EEEEE=7=?WanmcWOOYaYYROYgnngaaggnv�zwggWWRRO[\WOE<EOW\OTLA/)%-%-)..<BOTavvvnvvvvvva]jnaWaaWEABOTYaYOOE<<<,,),,-9BET]]Wbny��vvnOD<66/9=DObanv�����������������������������������������Ϸ�����������������ywpwv����z����zranp���wnmwzzwpa\aE6///5EYPEEOP\\amrmr�zzmrmrwmYYY\agmmhh\aagr�����������rrzaYPY\\mzrmaaYSJSYaSH=EEEJYJE=5EYgwwgROOYWWWYa\nrrwmaganz��yppgb[g[gnbOD<<<EOOWO=9/%%&).6BOTanav��vnvvaWTTLOWj]OLLTannWWOE<96/4//<<EBLOLLOWnp�vvnbOO<6649BWbnv�����������ż�������������������������¼�¼��������³���������zpppppwwvwvy��zwrz���z�wnnpnnaaYWR=6/6=HPYYYacamrmw�z�zwnahaa\\YYYaaamccchhmhwrrmzzz���rY\YH==HOYmwmaYca\YSY\HE=EJES\SHEEO\crwgaWWYYOY\\aawz��pgawz���ywpppppgggRD=<<<EEOEB6/,))).<BDLWbn����vnnabWWTOWWOELOWnnaabWO<6936<BDOOEEDL6OabnvvvannaO<<<=EOnn������������ϼ������������������������¹������������¼���������znngng\aagr�����z�����wrgnYaag\\OO=8==EYannwwrrz�����zwrcacYSY\\YYaaaghmhhhmaZaYammmrwhYH85/15=PYmnmaacmrg\SSOE==JSYY\OOOYhmmzzgWWaWOORWYgzz���www��������vvp[RROEO<<<<=EB</696*)%/.69EWan����vvnanaWWWTOEDOWbnbWbnbOE<93BBOaWWO<B96aabnnnnvvnaOODDEOap������������ϼ���������������������ѷ���������������¹��ż���znpnaWWWYYg����������wprrg\YaaYWO??EPPYczz�����������zzrha\YS\\\YY\mpzzz�zhggca\Y\PaaaEE6*!!$+8EYhhaYacr�raYPO?EEPaYaYSP\\ggmzzgYaYYEERRgpw���������z������znY[WRWWOE=<<<<=<<<6/.%%%%,)/<Tnvvv����vnbbWbaWYOOWWbnbWbaWO<<<BDOannnaW<4)nbnnnanv���vvnaWOWWn�������������ű�����������������������Ť���������������������ų�vy�nnWWYYYg���������zngnprngnYOOE?EP\\mz������������zz�zrha\\\S\\\gggz����zrg\\\\S?JPH5/*!$=Sa\Yachr�zmaWYPPYRaaaaaagmanmrpgaYOEEEYgzz���������www������yn\WOW[WE<766=ABA=66/)%&%%)6Oaann�����vnba]]aaaaWbWWnWOWWED<BBDWnvvvnna<6,nvvvnnp�����vnnbnp�������������ϼ���������������������ż����������������������Ҽ��zzznW[YW\w���������znannnnnn\JOYYEYam��������������z���{fg\gYRYYggmmwz���zrcYYSYE???81*	!2PSJPPchzzrha\acmaaanwmagmaaammaaYE=?EEPhw���������zrnwz�������vpaROWWE6<<6<B=<666/*,%%4BOOavv��vnWWT]annnvbaaWWOOD<6<LODWnpnnnaWD3%��������������vyy����������������¼�����������������ż����vv��������������������Ũ����znn\aar���������wnYS\gwng\\\naYacw��������ù����}��zrmccmcYY^clcmmw���xwmcZPF=/**++*=?JFESgmrmgaanwwwnnmmmrrngYYaaYYaO=5EESn����������wwpz���������paWHOO=.6<<6<=7466/%,6<DObnnbnnba]TWWYnvvnnaWWOOE6//6LDLTbnnvnaO<.������������Ż��������������������¼����������������������znvnv�������������������¼������wprrz�������zrnaWY\grnpngwrmamrwz����ý�ƾ������zmxmmchmhccZZhhZcox�{rsoeQA5*!*15=?P\hgnaaar�zzzmcanmwmaSOOEEY\J?=ES\p�����������wz����������vbWYH<6<66<46A<666/%%%,%.6<ETWOWbWa]TLTOnvvnnnnWOO<96<9<DO]kknnnWD9,�®�����Ż�����������������������ϼ���������������������vnnnnnn����������������Ƽ�������zzzwrw��z���wgaa\\ggngnwzz�zz������������ƽ�����mmcmsohfsf`XJXZXSXht{{sseX;1"$!$2EEJcmnaaar���zmaaarwmaHH=?<HYHEPa\ggz����������zw�������zvvgaYYH<6<<.666<6=</-/)%%-%%%%,,.6DETWOWOOOOWavvnnvaODD99<LE<BOWaknnbOD.%���˻���������Ż�����������������ż������������������vb[WWgnnnnv�������������������¼�������wrprzzppwpr\aYnhgg\w�z�����������������Ƴ����xhZes{trmshZXPPPPJJYms{rhZJ;'"&*!#++1?EYamcam{���wraPahmraOE8=8OPSSYhgprz�������������������zvnaaYWOD<</.6<64666,////-/%%).<DELOEEEObnnnnvaaOD<<99BEEDWWWabWOL<4,%�������������������Ż������������������������������vpWOLAO\nnvv��������������������ż��������zw�zrpgpgaa\nnmmngz�������������������Ʃ����sefss{{{wmcPSJJF=HEP\mmzmcP1$!--!!$$*8?PYahhmz����maSWchmYEE=7=EY\a\cmzz���������������������wa\WRODD<666666//-*4/69/)%)4<BD966<OWa�vnbOE9.//9<BEWbWakTDB6/%�������������������������������������ż�����������vnnWOLOOWaan����������������ż�������ż�����z�rpnaaaWaanggmnz��������������������ħ����ssrrr��{zrZPPPPF;=?JSamrrZP'""((&*/8=PYamm�����acYYc\\O7882=Raa\cmrz����������������wpwz���rbWOE<HE<<<666./)/46696/)%.66,%.9Lan�vbOD<6),49DOWbWTTDD<)%��������������������˱���������������·����������vnW]OETWYOYanv��������������±���������ű�����zg\aRRRY\ma\\amw�������������������н����rwrw{{��{rmZYPJ=5588FPYmmaY=*!!""(!$+6:=Pahm����wa\\a\YHE8525=Snaagzzw����������zw����wwmpzzpnYOEE=D<<<>6.).)/69==<9/)%%%,.,36DWbvvvnO946%,66<OWTLIB93)%��������������������������������������˼��������vbWWOEYaYYaav����������������������ƴ��������na\ROOOYanmaacgrz������������������ʽ�����{r{����wsh\Y;=555=88PPYYJ;1!!!!!$""+8?HSchw��zrr\\ZYPJ?=58?EPggrrwww������zzzzz������wnnpnaaaYWO=DD<D><,)).6<AEAA56/*)*%,,,66<OWWabaO63/%%,6/EEB<934%����������������������Ż���������������ŷ��������aWWTOOPaannv��������������������������������nWYYRWWYanrrggcmw�������ƾ���������Ľ���z�{{�����mhYYP8++15==8?FF?881***!*!$$8ESZ\hmrmhmZSJJPJE=?E?ES\rzzwz����zwpwwwww�zzvzrnhg\YWaYaaWOEGODE<4..6<DLOOOEEE9//*/-%%%3.36DDDOWD9.)%%),6<B<6.%��������������������Ż��ų�������������¼��������nW]WROYnnnv���yzzy�z��zppvnnz���������������wn\YSYWRanngrmmhz�������ƽ��������ư����z{zw����zcPPJ=1*+1855===?8581**/*!!18JS\ZSYYZZZPEEFJJJJHHSYYh������zrmaapwrgnzrrnngcWWOEOOWYanWOWWOE<<63<DORaaWOO^TE==/*-%,.333,69DOD6%%-,%)%/6664/%��������������������ջ��ż���������������������vanndngnnvvvw����rnnnvgnbWHHRHRgwvzz��pzw������zgWYYYO[gwwrhamnz�����������������������rhmm��{rhZJ8511**'18111111+11*'''!!&18?SHFEFJSYJF=?JJJPScc\Yr�����zwrraaggmaaaa\Y\SOOO?<E?EPYaWYWOOH>>><<HRa[\YWO^aOOL/)-&)%)43)%.6<B9%,,)%))494/,%���������������������ϻ��Ź����������������������vnvnvnv�������wnkaaYOD><66/=Wagannnarr�������gWaYRamwzzwmgrrrzz������������������zwwmcm{�{r\aS?5/'*++1151''$*$$+11551*+!*58?J=11=JYFE=?FJPYhmhcawz�z�z�zraYYYY\\PPYYPEEE<66666EEOEPRWOHWOOOEOR\npnaaaWTWWL=*)%*%)%))%,334)/,%).44,))%��������������������������ϼ����������������������vy����������vnkaYWO<<.)%%/=OWOOW\aanww�����rnnagwz�zzrrwwznnw������������mmmarmmmmcYm{{raYSJF1+$*''1151'$!!$1=?=111*!"-5188+*5;?HE=8=FSYrgmhmz�zwwz��mYHEEEJYOO?==<76+!%*4=?7=EOOWWWWWWWaanpvnaWOOEEL9//**%,,%%%,/,)%,/-)%

����������������������������¼�����������®��������������������pnaaO<6///=E???OOWgp�����zrvz�������zwzrwhapz����������cSPJPSYhmmZPcwshYSJ?;5'"$$'58''$$$!$108=85+**$(511+*'18=?=88FScrmmmmrrwwww�rgSEEEEHOOEE=62**//22EEOWRRRWWbaaanwa\WYOEE<96/*%,,)/64.))-.-�����������������������������ż����������¨��������������������wnYTOO=/+#+7866/7=P\r����zprz�����������rmahm���������zrP=8558HYcZZZcmcZP;;81($$$!'01'*$"!$+188+1'1'$$"1*!*#$*/58858FYcmnaamwrrrwzwra\HHHPEFPE=772**/66<EHHHHOWWWWWWn\WWYOE<69<6%,,
),6<9,.//.������������������������������ű�������������������������������nYOTOL6**68<*)+//<Jhz����zw�������������wwm{���������rcP5'***8JPXZcZcZPF85'*!$$'1''$"+11''1111++'("("!!!#+**'15=FPYaaYacmmmgmwrga\WWYOYSSO=<6/!#*68=HHEEHEOEE=ERWRWOL96966.%%%)%
)%,..,./3/������������������������������ϼ������������������������������zaOOTLO<#)/7/##+6??\w�����z����������������wx{{���w��zmP8'$!*1;PYYYYPJ;1"$$+11+$$$$''11811081++$""""#+$**15==EJHSaaaammrrmcagaSYYa\PE?=/#*/7===E96<6<6<DOOOB6///6/%))/..,%%%)%%).4/..�������������������������������ˮ�����������������������������zaEOOLE6.)*#+/664*))9EYagmrz�zz���������������wmrs�{�rmw��cP=+$1;SZYYJE;1*$11''"'11888;;81'!$$!**'''"!$+!!**1155EJYaaaawrmhgcrga\aYSSOE?/
#/2786/*).+/6<<6<-**%))%)%,<<96,.,
-/3,%
����������ż�������������������˹�����������������������������rkOOOOE>66//626<<=676++9ES\YaYcnrwzz��������������{s{r{��www�wmJ5$$2=FZZYF81($$!*''''''0;;JNPJ;8'$$$*'!$*'111!&&*++*!!!*(5=ShnaaamrrrrmmhaYYPYYP?6*#)*)***%#).6/),,),3<DEL<3.)%%-�������������������������������ϼ����������������������yvv��wwaTWYRO?>6<DWE=EEH=E7<<=S\ggYWOYnmzzz�������������{{{z����xrrmZF5+*!*188;PZ\J8$'''0'1''''';NZZ`XNJ1'$$'1''1118;1'""(-1++!!*8EchaaccwwwmchaYYSPSYPE6*!)))).)*-.9DOLIO<<,/))
%����������������»��������������ϼ���������������������nnnnywnYWWWOHODDDHWgWRWYOOOO?HP\aaaWEOOWhnzz��������������������rmrhaYF=55/*5;=FS\X?1'18;;0''+'  ';Nhhr``XS8''"$''18;5;;?881'11558/!!1?SacYYcrmgcZYSYYRYYYYE=+!)-49DOOOIIB6<4/,%�������ű�����������������������ż��������������������pnannnnWOEOTOEDHRWYnvpgp\REOWaa\gaaaYOEEEY\mwwrwrw�������������zrwmhYYPFF=8558F;JJSJ1'" 0;;?;0'''             ';N`r{ttrhS;8181'18;8;;?=F;;;;F;81**18EJOammca\ZYOPHSRSOOYPE2****4<DOOIDOB6D<3%.�����������������������¹�����ż��������������������vnnWaYWYYOE9AOHEHOabnpy�vnOOWkwwvrnYYOE?8=EY\ahhnrz�������������{{rmcSYPPJJ????F;FSJ?0'*'?SNJ;0' ''              :;Zs{{{{f`XS;:80;8?JJ;;?EPJNKFF;82$*11=;JamacchYOE8=EJHYYPE?6*
-///6ABDOODDB7<<3%.�����������������������������Ů�������������������vvaWYWWLOOO<<6DHHERWYnpz���raYWgr��zznWO=6?EPYYYSYarrz�������������smYZSPJPPP;JJF?;SSP;81'$'+8JXV@;''+''   '  '       ':N`ft{rff`hXJ;;;;;XS;JPJJXhZZQF;?2$$*15=JYY\YaaYE=58EHHOPE</*


*6/46566<OIOD666.%,��������������������������������������������������vnnkYYOOLAEEEA<DHHHRRb\nv��wwWOYnw����zcY=28?EOEHHSarz�w|{}��������{rZPJFPJJJJ;;JFJ;JJSJ;;01+ ':;NXX;00''0000'0''        '0;NXffhsff``ZVNNNXZSSSSSSZhsfcPP?7+!**115?PPYaSPYP?516===EE8*
*//6666DOOOD<6.)

%/������������������������������������������������vnnnnnaWOE<EOEEEEHHOW\[pvvvrnYOYw������nYE56<=EEESSarz{xx{���������whYSF=FJJ?FJSEFPJ;SSS;;0800;;N`Z`N;0000;;;;;;0'        '0;Nff`fftsrff`X`hXNSXSYShrs{shYP?:15588;FHSYSPEE=5//22////*	
%*/4444<DIO<B/,)
%./6���������������v����v��vvv�������������ynannnnaYWOEOLEHHOOHWW\WganaaaOESnz����znYH==58=EJHYpprmso{z�������wrcZSJEFPJFJSJPJP;;NSSSJCJNNNXZ_``X@;00;@NNNN;;0    '   000@Xffff{{t{t``fhSNSJSScfr�{{soxcVHJJJ?;J;PHEE=11**!*$$!!	#*+
)///6LL<<3,%)/6<B9����������ű�����yvvanaWanWWWanvnn�����������vnkknnnvnnaWHEBEROWRRWW\WaYaWYEE?Hg�����zvYOE=78=ES\gprmccorzrrmz{zwmmYYSYF;?PSSZXSSPJJ;SXXSSX`hf``fff`X;00;@XNX;;;00' 00   000;NZfit}���}t}{fh\SVVhhrr{{{�����rrhZP;FF?O?=//!						)+/+%/4==9.)



/9<ABE94���������ϻ�����y��vnaOE<<BE<9BLTOTWn���������vnnnkavvyynWE<6<HRWWWRbagWYYYWO>6=Hg�����znaSE6258ESanrrnhhemrrhammmmmhYS\ZYFHJPZZZSJJSSSJXXVhrttifitff`X@;;:;@@@@0;;000000000000;N`t���������tthZhZhfrrst���������hZJ=EF?8(*$								$*!)/2/+)44,)
%%)/69IB</%���������Ż����ypn�vnaOA66,...669EIIOWn���vnnnakknpaO>66<<HOW\\a\WYOOYaO<6=E\����zvg\\O82*5?Pagmmmmha\h\YZYccZccZccYZSJJSSZZZJNXSSKS``ttt}tt}qtf`X@@@@@@@;@;;;000;@@@;;;:;;N`f}��������{tffh`r{rhrr{���������oP==88'*!				!*)///+))&
,4)%)%%,.,6<<D9))��������������nnvvbWB46)%%..6BOODOWa�vvnvnnaaaaknvpnOE966<DDEEWaWOHHHHOaOE=EEYarzzzra\\PE=//=H\hmhhhZYSYSPYPZYYYZ\YZY\SJJJSZZZNSVZZXXfrft}}}qttifXXXXVXXXNN@N@@;;@NNNN@@@@;;;Vfq�������}�{ts`hftrhrr{��������{hSP?5*!!						!!!%/////6/*))#)))%6664.,,%-,6/66<D<</)v�������������vnvnnTE6/.%)39<DDDOOWnnvvngnnnnanank^YE6/6<<EEEHRWWE??HEW\WHHOHRYarwwrnaYPPE828ERammcc\SJPPHJJYYSJPSS\\ZSJSSSZZZXVZ`XVX`ftt�}}}qiiifiiiiffffVV@NN@NffffXXXN@@@@Nf}��������}{trffhfhZr����������trYJF'!							*!!/666/66/)))%,3<<66,),)669436<<66<<66.)nn����������vnnnWE6,).6B<DDDDOOWavngggnnnnaYYPEA<4466EEOEEHWWOWOOOWaY\Y\\YY\gmaaa\\YHE=8<>P^ceoZYSSF?888;JF?;JPchmZSXZZhZZZZhZXNNXfq}����}qtiffiiffXfXXNNNNViq}}qiiifNXN@ft}��������}{fhhhhh`hz�����������mP;5*!								!!*)+//+/)*,69<3,,%//69B<<EODE<B44.6/nnvvvpnvv���yvbaLB4,,<LIEOTOODDOa[[YnnnaYaTPE6664466<<E<6<=Ra\YYaaaknmpnmaa\YYYgghaSHEE>?HYZZZZZ\SP==585=588?S\hhZZ\rs{trhZhZX;NVft}�����}tiffifi`VVXXN@NNfq}����qqiifXftq��������}qf`VVX`hfft����������zhS;1*								)**))*)/696.,%%.69<<<BEOODD9,%%,)nnvnnnb]bWnv���yzbD64,,6DEWOTIID<<EORS\nnaYYaTL6/,/6466.<E<66=R\aa\grzzr���raWWWOYamnYSJOOH?EPXKJYSSPF?=8551118;SZhhZZh{{}trf`f`N;;V`}}�����}}ifffiffNNNNNNNffq}������~}iiq����������}tfXXNNVttt}����������r\?=1$								!!+
).6<6,%,3<66<BOWOEE<)%%annWWOODLDWnv�y�vaE/-%%,6=WWW]]OEE<EOIOannnaaaYE6*%%-//)/<EE6/7Hagnmp�������wgWWYYYS\aYSSOOHEMSKJFPEE=;=;55515125XZh`Zhs�{t{tff`Z;;0NXt}������}qffitifN@@@NNfiq}}��������}}�����������}qfXXN``fttt���{{{���xcN?//!					!**)	)%336,%%%.<<<6<9ObWOOB/aWOOE<936BOavpnOE4.)%%6<OWbObkTOB<<DDEannnpnnaE4)%)/666<<</6<EYgnnz��������naa\YYJOYYSPHNEEFJ;;EE?8515F=5111215FZhehf{{{tttf`VN;;;N_ft{�����}qiiqqqiXNN@Niiqq}�����������������}}��}}ifXXN``fsttt}{rhss{shP?7*!!		!!!$**//!%,.36,%%36<<<B9EWOWOB9/bWOE<B96<DWavnvpnnWB9,.,.3,46AOWbbbnb]OB6<DDESnnvvpvkE6/))-<=E><<6/6=H\pz����������p\\\YPHHSYYHHH=FFK;?==?5515585858118ESZZmsr�{tttf`X;;@NV``ftt}}}}qtqiqqqqifffiqqq}}����������������}iqq}tffXNN@X``ssttttrrrh`XF;12*!$$/+*$$**/1*

)%,)694)%.36<<<BLLWWWD64-,%aWE6<399BIObnnvyvvWOB3..666<OTWaWbWWWbWOBBDOOgnvyyynYA644<<D??E<6<<=Rp������������wgYPOPPPEJOORHEFFK;====888=;5858=11=?PZZhst{}tfff`N@@NVXXfifiqtqqqiiqqqqqqqq~~~~~~�����������������qqqqqifXXNNNXX`fsfrhfrfhSSK;5++$!*!**$/62/$*/*+*


)%)%)%,669664,499BELTW]OB4--/naO9639BBDOOWnp��vTTL<<<<<EOaaWaWOOOWWOI<<IOgnvv��ypkOE6<OE=EE>>DOOOay�������������waYPOHEEEEOSSMPK;?=8=?FPJFF;88;;;;=FJSZhrt{{ttff`XNNVVXfttiiqqqqiqqqqqq~~~~~~~~~�����������������~qqiiiiffXNNXXXXX`XV`hfZVJ;;11-$!$$!*+/$$+///*//*!)#)))%%,,,,%%%449<EA<4..699ELLEOE94)%vaD996<<<<=<Oan��vbWOOEDLOOavaaWOOWWOTTD39DYavy��vvyvnYOOYWDDDDDDWWWn������w�������zn\PE===E=RW\UP;;5588=ESSPP?;8;JSJJJJSShrt}�}tf`X`Vfff`ittiiqqqqiqq}~~~~~~~�~�~~~����������������}qqiiiiifXXXXXXNNN;;;SXNN?8'01($!!!*****!$$$+66/)%))6.)%%4.66<36669<LWTA4)/6666<<6/%vaOE<BBBB<E<OWp��vnnnaWOWavvnaYOOWWWOD<99BOWnv���nv�naYgWRE><DOR[nn�����zr������znaYJH===HHHSYYP;85/188?JYYSPJFPSZ\SZJNSZ`htt}}ff`ffft}}}}}qiiqqqq}���~���������������������������~}qiffiiiff`XNNNN;000;NN;81'''11$$*!!//2/*%
)/./6./,-%%636<D<<<69LYYYB6%%,%),43)
vbWLBEILEDOOOay��������v�vvnnkOOOOOIB99D<DOYnnvzvyy�z�nnaWOEDDWbgvvv����wrwzzrwzvg\OEH===HEHSYPF;55/588=E?JJSSSXcmhhcZSSSVZ`fftfttft{�����}}iiiqqq~��������������������������������~qifffifiifXX@@;0' 0;;;?01''11-$		!*+****!
))666<4//,))**46-%,/6<IWOD<<BWWbWE6%%)%,%
nbWaTTLEWWWWWv�������������vnbkWO>DEO<6<IDEOWnanv�vvpz����ga[WODDOanyvpzw�znaagg\mnnaSEE=76==?HHUP;E58888E==FFPSZZccrrrhZXSS`ZVVX`tq}{}�����}}}qqiiq~���������������������������������~}qqqiiiiiXXX@;00 '0::001'+"''1$						!**))!*%#*%)6<6<AB6/6//6<<=96669IWWWOE<LaanbE6)%%)nabnn]WWnnnnnv������ű�����nnbWDD<<<<6BOIEOYWYanvnnnw����znabWDDOavzvnannwYOORSR\\aYJE788668?HPYS;F58EFFPJYPPPZZZccrx{hhX\Z`VN@NXft}��������}qqiiq~~�~�������������������������������~~~}qqiiifNN@;000'''+''1'''1($$!					*66/*-**//)//66/))*)))+/6<?OOB<A<==LYYTOOE6<OTbajTT]WnaW9,))%).nnnnvpnvnnnv����������˼����nbOEH<<<DDOIAEOEOPakaaaz�����vpaWGEOWnvna^aknO>HEHOOEEEE62/<==ERSPPKJE=FPPY\hhhh\chchhmz{rhZ`ZVNNNNVftt���������~qqq~~~������������������������������~������qqifXN@@::00+''   ' $'"(*+++$!!							+==6/*#-/+/6466<7<666/666.6<HRYWE<=OOOYnannaOBBObnpnbbYanbO6.,,)))%vnvnvv���vvn�����������ռ���vbWEHDEDIORDLELEEOYYYYYw������pgROEOWgaaWOOOOO??E?E==5==2+/5?P\_aYPJJEEPYYZcmmmmrhmhmhhszrshrfVN;NVff`t����������q~~��~����������������������������~~~~~����qqqfN@@@;00' +'    ""111'*					/266//**////6>?H=<<E<<69<<?>EWWbWOLLOYnanvnpn\DOYnvynnabaWW<63,.)-bnnvnyyv�������������ټ����vnWOOOWODDIOOOTOEOLOYLYn������ppbWWWWgaYOE>EE<7<7<=2266565=7=YgrmcYXSEJFYY\cmmchhrmmmhh{{tffsf`VNNXfft������Ķ����~���~��������������ǿ�������������~~~�����qqqfNNN@;000       "('0+**$!					&*+52/*-//76?OROOO\\OOOHHOOOWORY[\^Wnn���yndWbnvnyvnnvnaWWO<6/),bnnvppv�����������������ż���nWYOOWOOOW[\aYWOE9AELYaw���zzyvvnnabaaYO<7?<=666622+/665=E=OYgpacZXSHPPPSSY\YYYZhrmhhh{�{trrf`XXX_ft}�����������������������������������ǿ���������~~~�����~qqiffN@@000'0'    !$++$*!!!!			&//52/667<6?OaaY\vpnWa[aROOOEEHRaap��������vvnnvnnvyyvnnbbOB<.%,an��������������������ϼ±��vnYYYaYWWana\YOE=<AOLYYn�������zzvpnnaW?7666466/76//6665=ESO\grmhZXPEYPPPYYYYJPZhw{rhmr{}{rtf`XX`itt������������������������������������ǿ���������~~������~qiiiifN@@0000'        !+ $!!!!****!								/625<<6<?<?Okngry�yvnnpgWOOEOOR[w�����������yvja]nn���yvvnnbOL9)
6nv����������������������¼����naaYannnnannnY?=<6EOPYYa�������yzzvznWE6//.*///*/2+/=E?=EJRSY\nwmZXPJSJYPSZYXSZZhw{xrrrrt{�t{th`f}t�������������������������������������ǿ�����������������~~qiiiiNN@@0000      $$$!!!$'+*1*!							!68EEE<==OYnwpw��yvvpvaHDOWOYgz�����������pn]ann����vnnnkW<6%,6nv������������������ż��������vnnaannnngvpnaH?=BOSYagn��y���zyzzvynO>/)*)*+/*/266?POYSSSSY\nwcZZYPSPSPEEPSZccmw�{rrrfrt}��}tft}}��������������������������������������ǿ��ǿ�������������~qqqiiiNN@@;00     ! !$*1'11((*$					*5=EOE=<HYmrzw�����yzvpgRO<OOWn�z�����������vpaajn������vnaaE</)))/<vv��������������������������vvvvnavvgnnnaEE<AOaanwnnvnvvv�����naE//))%***)66??EYchaaagrrmcZZYSSOOH?;FYYchr{�{tsffrt}}�}}}�����������~�����������������������������ǿ���ǿ�����������~~~qqqqiffNN@;0      #!*1*11555=5**!				$6E?EEE?Wgnwz�z�����zbaaO<<EOWgwyvv��������vnnjaavv��vaWOE6464/)),/46vn��������������������������zzyvnvnngna^YOWOYapwpYnnnnvy����p\H<6/**!**/7OOOYamrz�rzwmZZZYSSH=8==FJccmr��{�ssrtt�}}}������������}}�������������������������������������ǿ��������~~~~qqqqqifN@0         $*/158?EHJ==/+!					+?E=<ER\gnnpzz����vWROD<<<EWYnpnnnn����vnaaWWbanvv���vkaOE<EBE9<6.4.4v�v���������vv�����������ynvnvngggnnaaYaWYYnznWWYbgpnz���pYE<62/!*-/=PPPYmr���rfmmhehYSS?=8=;FS\hrr{��{tttt{}}}����������}qqqq��������������������������������������Ƕ�������~~~~q}�qqff@;00'''    !$/5=HSSaYS=11**!*							5EEEEOWWgkwzzy��w�nWHE</9<<=OYnaaOYnvnngvvnbWOOOOWbnv����vnbWEOTTOED<99.3vvv������z�vvnnnn������������ynnbWYb[nnnakanaaWapWOHOWaWgv��vnYE=6/#*-/=EYamzz���zgmmsxshcSE?===FPZhr{{{{{ttrr`frt����������}qii~��������������������������������������ǫ��������~~���}qifNN@000''    $+88;PPYacYF5+*!**					/=EE<?RY\aaz�wpzvnaWHD</,/66EOOTOOOEEPTYavgWOBBDOObnv��vnTWWWbWOOOOE<9.nvvvv�����vyvnnanvvv������������vnbOOWagaYYWT^anYOYYH?E>OWWgavng\YE=7+)%!*****2?Ymrzzz�zrgmw{{xrhSYPHFFJYhrz�{s{{{rh```ht����������}qqq~�������������������������������������ǿ������~���~�~}qiifX@@000      $$+18;EYZcaYS=/**$!			*6<776?EEEYagYapn\OHED<./466/69699=/)/4EYd[O<<46EOWbabaannaWannvaWbWWEO<9nnnnv�����ynabbn���������������bOLW[OPOLLOYWnaWOEE9666OWWWWROOHE</6/+!)//**+2=P\hmmwzrgnmx���whaccYXXcs������{tshZX`Z`f}��������qqqqq~������������������������������������ǿ����������~~~~qqiNN@@000   '    ''"**+ $1/5=ES\SYJJA5/*!/2//6<E<E?OO?EYWWE<DEE6666./%%)-,%%4=<O<6646<DEEOEOOWbaWnvvnnabbaWODEWWWbnv���nnaav����������������aOOOWOEEEOOOWYWWO<6.)).<<EEGE?===7666//*/72/**/=EH\mmrnhggmw����xhhmcZos{�����{{tr`ZSV`fft}�����}tiqq}~������������������������������������ǿ��������~���~~~qifN@@00000 000++'''80'-'0+"'158;;JPPHFF=5/*$!!*+-//6<<6666//=EOE/<E><6.))%,36,,%/66<499<<OTWWnnvnvbnabWODEDWav�������vnn������®���������aOILII==AWWWWWOOB6/%)./66<=66//66=646726////58=5Pamgh\gpw������wxx��z{������{hhhhh```fit�����}tiiqqq~�����������������������������������ǿ����������~�~~~~qN@@@@00000 00:::0;:;;;5108888;FFF?JJE?=5/**+/*!!%**)$)-*//+))/)*/===6/66/),/.,%%,6<DOWWvyvvvnbppnnn6<OWav���������vv�����������������vaOOIDD=<LOWTWOLB6/))/666/)/6796=?7-////6676=HY\ggpz������������������{shhhrsshhft}}����}tqqqqq}�������ǿ���������������������������ǿ���������~~~~q~~q@@@@@00000000:;;;NSNNSP;:HJ?;FFFFE==855//*$$/6=76+/*#+/*$!*/66)))))
%%%%,39OWWvvvvvvnnppn/<Eav���������vv���������������vnaWLLLE=LOTOYWL64)/76+*)2?=>=<E=6////+*2676=HS\h�������������������shhrrr{rsst}tt����}ttqq}}~����������ǿ�������������������������ǿ������~~~~~~qq~qfN@@@@0@@@:;;:;NV\hZXXZPCSJJ8=FFFE85*'//*+*$**2EYYE==/+*/*)+)
%6<OWnnzvvvpnv��%6On����������v����������������vvaOOOEEOOLOOO<<%)/2226<<>E=???=7///**6226=ESnz������������������rhhrrs{{�}�{}}q}��}ttqq}}����������ǿ�������������������������ǿ�����~��~~~~qiq~~ff@@@@@@X@;0;;@N``fffsohVSSFF;?;;=5'!"*/*/1**2=SagSYE=6*!
)6<Oavzvv�yp��-6On�����Ż���yv�����������������vaWWOOEOWLTEA<<*+67=<6=?EHEE<222**+2656=APgv{�����������������rhhhrzrr��}ttt}}}}}ttqq}������������ǿ������������������������Կ�����~~~~~~~qiq~~iiffNNNNXN@;;@NX`frt{{xsh\ZXSPE;5/1*('1//161+<S\aaYSPF=+	
,49<Oy����vv��6<Onv������®���������������������vbOWEOPaOOB966)*/266/==?HEE767=2/++/6===?\pm�{���������������{rt{t{{����t}q}�zz�}}}}���������������������������������������Կ������~~~~~~qiq~~qqqqifffffXNNN``ftt}���{rhc\XYPJ811515555==8=PYaa\YPOO=/!,4DOnv�����vv�OOWnv��������¨��������������v������pWOYYanaO96/6/)-%))/**/66<<<<<<E=?62//6/62ERghws{������������������{{������}}}������������������������������������������������ǿ��������~~~qiq~~}~~}qqqtttf`````fs{}����zhhZSZYS?8=585=FPJJFPPYYY\aYSOE2*
3EObbn�������Wnnvv��������Ź�����������ypnvv�����nbbaanaWE=///<=6,%#*)///2667EEE?=56*6//5EW_ruher��������������{��������������������������������������������������������������ǿ�������~~~qi~~~}�������qqif````Xhtt{���}xmcSSSJ;=8=5==J\\SSSOPHHSSPOE82*



)6BTaa��������v����������ż���������nabnnnnnv�ynnpnYaaWO=<647HH96))++)*)%#%)*+//2EROO?=56**/=OS\\ccXhw�����������������������������������������������������������������������������ǿ�������~~qq~������������}i`ffZVhrft�����whYSJ==8=EJEES\ma\YEOHEHE=E56*


%.9<Wnv������������������������ų����zvaWb]bWabnvvnpznaYOOOEA<==OOEB<6/6/4/2/**//<EWRRJE?2*$/=O\\\aYXXh������������������������������������������������������������������������������ǿ���~~~~~~~~�������������}tff`XXhet{�����mcS;515=PSYZcmmma\O?EE=76/2*!)%.9Obv�������v����������������ŷ�����vpnWWbWbWWaannnp�zvaOOWOAA===EEDOEDE<<6676+**/<HYYSPP?=/++/?H\SaYZZcm�����������������������������������������������������������������������������ǿ����~~~~~~����������������}rZ`Zhfs{�����mcSF5/5FPYhrzzzwcaEE=/6+*&*!#.)),/)6Dbn�����n����������������ų����vpaWWDOWWWanvnbnpvnaaWOE=66==EOOOHOOE</62/)*=S\\aYYFE=7666H\\achhmhm{w�������������ĵ�����������������������������������������������������������ǫ����~~~~q~�����������������thhhhtt����{zwrcJ;1=PYmw����wmcS?2+***)$&.6/)//,.6On������nŻ��������������ż������vnWOEEOWnnbnanvvvnvnnWE<=4<EOWYWWWWOE662/-**6EWanaaYYPEEE66P_gnwxswwwrww�������������Ľ����������������Ͷ���������������������������������������Կ����~~~~q~�������������������{rrr}�{{{��wzwhYF;EScw�������mYJ6+$***+6366..
)3<Wv�����n�����������������˼����vaWOWWbnvnbnvvvnnWEE<6EOaWggbWOED<726/)#*2=OYanvaa\OEEE=EOgz��������{���������������θ��������������������������������������������������������ǿ����~~~qqq~���}~������������}{ttt}��{}t{rrraSPPPSmw�������rhS=2**/*)!*-	)6/.66/#
%),9Dnv����yn�������������������Ů���naanvvvy�vnnv���v��nnYOL=AEEOW[bkW<6<E==676///))*/<OYYYannn\PE=EHS\r����������{z����������������������������������������������������������������������Կ�����~~~qqq~~~qqq������������tttt}t{{�}rsrrrYSPPYYcww�������raYE8===5/+/**/*).)/6),)).3DWn�����n�������������������ձ���nv����y�y�������vnaaYAOOOEEER^aO</6<=E<E7<76///=HSYYYnnraYJEEHYarz�������������������������������ĸ�����������Ͳ������������������������������������Ϳ����~~~~qqq~~qiiqq}���������}{trt}}{{ztrrrrrmcSPSYcm��������zrnaPE?FE?88<72/)%


%).<<Oav����v��ŷ����������������ű���������������������vnaaTLEYA<>EOTWO<./6EOEOOE?7/66OYaaYanaaa\YEHYagw������ʽ�������������������������������������ʶ�����������������������������������ǿ�����~~~qqqq~~f@ffiiq}�������}{}}}}��{tt{rz�{{r\YYZcrz����������raYOYSPWEOE7*	
%%%%4<DOapy�����������������������Ϸ���������������������vnaTOAALE<<EBLOE<666=EOWOE?=6<=OYnnYYn\Y\hYYYYam���������ƹ���������������������������ĭ�������Ͷ���������������������������������ǿ������~~~qiiq~i@@@NNfitq}�������������{}tsr������rrmmmw�zzwz�����whgn\ggnaYH7/
)))

,4<OOWpy��ű������������������ż��������ż�����Ź����vaE5=9<<<7<EDEO><<E=EOOYRE?=?HWgwraYYW[\aaagarr�����������ƽ�������������������������������������������������������������������ǿ����������~qqq~qf@@@@Nffiit}}������������}rsrz�������xrmhcaawz�����wz�zvwz�waOE<*
))#)/+
)6<DObv����������������������Ź����������������Ů����vYA=666<<EE=DOOHEHHD=OWa\^POHRap�waWWWa\a\mmz��������������ð�����������������������������������������������������������������ǿ�����������~qq~~q@@@@@@NXffttttt{}��������}rmrz{�������wwcSYYnz���������z����wRE>2))/)

%4<BObv������������������¹��������������������˳��vnUE666E<EOEEAWaWWRWHOOYnga^YW\m�zn\RWY\\mrhw����������������ú���������������Ľ�������������Ķ����Ͷ��������������������������ǿ�����������~~~~~i@@@@@@@X`ffttttt}���������{r{zz��������whYPYnzz�������zz����zgS?7*))*)).<DWnv���������������������������������ϼ��¼¼���naL=666EOLOEEOYaa[[\RWWWnnvaampppnaYYSYR\anrz����������������ѽ������������������������������������������������������ǿ�ǿ�����ǿ�������������~~qf@@@fNNNNXfftttt}�����������{w{�������zzwmgamammwz���zzwnz���znWH</+)#

)6<<DL]nnv�������������������������������ų����������vgOE596=<EEEEEWYanpg[aaag\anww�pn\\OSYSSYJYmw�������������Ľ����ƽ����������������������������������������������������ǿ�����ǿ�����������������~qiiffifNN@Xffftt}�������������{{�����{���rwmraaYannmwrwr\\awz��pYH<644

,<LDOOTbnn����������������������������¹������������v\L=A=6<<=ELOTaanppnnnnngYYkw�zwYEE?PSPOOEYp���������������������ƽ���������������������������������������������������ǫ�����Ƕ������������~�����~}}qqqffXXfiift}�������������������������rzwwn\HYSPHYahYPPO\gnnaYO<<<<4/ALOWTTOWnn��������������zyyvpv����������������������\E569E66<EOaknnnnpnvparngannwzgWE<<?HEEERn����������������������ĽĽ�����������������������ʸ�������������������������������������������������������}}iifitqift���������������������z����zrwwm\HEOOEEOOE?===OWROYOE?E?6)))%6<OOOWIEEOO�������������ynanb]bn�������������v�������v\LE=EEE6<EYkvwpagpnrnaa\\aanmnaO<66<<DEO\n���������nrfmw{��������ƽ���������{{t������������ĸ�����������������������������ǿ��������������������������}}}}q}}�}��������������������zwr���rr{wrhYSPE=EE?55/6/2E?OHOEE?=76*)/),4,%%,).6<EOTOOOL<9<������������aWWWOT]avv����������v������v\OLOOWOOLTWavvvvnwgng\WR\gaaggnWE7<<<<OYgp����ƹ��zm\\SZmx����������������{mrss�������������������������������������������Ƕ���������������������������}}�������������������������{xmrrzzzzwwwwmhYPEEJ?=5/*)/77EOYP?E?==6-*%*/,),4.)%%6<BDOWW]OOOD</,�����������nWOOOEDObav�������v���y�������vaY]nnaannaaganngnn[RRROW\namnnaYH<>OEOW\nz����ƺ��wmSPRScms���������������smZhs�����������������������������������������������������������������������������������������������������mahwzr����zrmaSEJHE62/*6<==EE?EEEE</2*



/-/.,,4.,%%%,,4<OOWbbnnWWOE9)����������naWODBBDIOWv�����������������vnnp�vnw�znYYaaWRWWWOHHOWWYaaana\YOHRRR\az�����é��wcYEHHPcms�������������{rrhst�����������������������������������������������������������������������}�����������������������������wmmrrm����zrnaSHEFE=2/***/2=??OEPOEEE77+*44,),,.,%%%)..366<EWWannnbWOD63)����������vnnWO<.BLOObv�v��vy��������������v����vvnaaaaOEOOWODEOWOW\Ya^aaagna\Wgz�����Ƽ���mYJ???Hccm{������������{rmrr����������������������������������������������Ͷ������������������������}������������������������������wwzmmrzzzrhmnYHEOE888/////<<<EOYY^YOE</%#
%,.%,,,)%%),6BDOBLOankabWTO<6,),����������vnbOE9.<OWbbnv���vy����������������������vpaaWWOEOOODD<DEOOOYSWaamgnpmrw�����Ƽ����nSE==?Sammfs������������wmt{������������������������������������������������������������������������}���������������������������������zrrmrganrwmYPPPEEE=<=<5==EOYaanaYWE64%).6.)%%%)%%,6BLOOWTWab]WOLED<6664����������vnaWD99<ITnkvv����������������������������pnaYHHOWOE<<D<=EO?=?Eanwpwrz�������������aSE=8ES\mm{{������������{{{��������������������������������������������������������������������������}��������������������������������zwrragrz��zmcaPPYWOEEE?=ES\\gnwpnWO?</+)6<<6%%%%6BLWOWbjabWWD<<<<<43<9�������vnbWDBB<DTkny�������¼��������������������paYOELEEE<6<67=E<<7Ogzzz�vz������������wnaSWOPS\a{�����������������������������������������������������������������������������������������������������������������������������zrmrhr�����wm\ang\WRRRHHS\nrggnnaYOO<D<6)3<D<6)%%%%,))<OWWOaabYWa]O<A9E6699E����vnnnnaODBLEOWvz���������������¨�v������±����zaWOEB<<<66<6677<EOYgz��zzz�����������zmrhgna\\grxx���{�����zrw������������������������������������������������������������������������������������������������������������������zwww�z����zzzzzrpggYaOOawwnmmrmnYWWWOE<OOWHB4%%,%%,,.,,DWWjnnnaTWa]WDDB<<<<DO�����vnbWaanbWWOTTbny���������������Ѽ���������Ѽ����yaYHEE<66./<7666=OWamv������������zzzzzzr���zrrrrrwx{��zwmzrrrz��������������������ĵ��������������������������������������������������������������������������������������ó����zzw��wz����������znna\anwwppnpnngannnWR[an\W<6//.))%%%%6BObnpabW]WWTOEEEB<<EOW�����vaOOOWnbnnW]npv����������������Ů����������±���ynaYH<666266=646EOanvzz�����������vncmwz�����zrrgphwxs{rmmhrrw��������������������ĸ�������������������������������������������������������������������������������zz�������æ����zwwwmr�����������wwnnnnrwwpnaWagpwwnvnnp�znW=66-))).4,.9DOnvvabYOEBBDEAEBEDWb������vOOOObnnnaan�zz��������������ű����������ŷ�����vwaWE6/7=<E<462EOnrvvvwz���������nacmwzzz���rgma\\cmmoohchhmz����������������������������������������������������������������������������������������������������{ws�������ó������zwmr������������zz�zwzwvvnaW\gz��z���z��vaYE6///%%)3/.469BDWnnbOOL<9<9<<LTWbnn������nbWOWbnbannpz���z�v���������·��������������������nWE566<EOH==EOYnpnvnnn�������zrm\armwrrz�zrh\\\\YZ^ZZhZZhhz����������������������������������������������������������������������������������������������������{{�����������������zrz�����������������zzyvpaWav����������wnYOE=EA4%%),4496EBB<O]nWOB<9969<<Wnvnnv����vnnbbaaabapy�����py������������������������������nWE<666OYYHR\Wbapvraan�������zwghmhcaamrmnnaaYYP\YUPXZSPXZz�����������������������������������������������������������������������������Ľ������������������������������������������w�������������������yngYp������������vwnaWOLB-%,,36<B<ELLEEODOE944/99<<Tnvv����vnnabnaabbv�������zy������������������������������nT<9<6=EWggnnggv�vrnr��������zwrwmnaYagna\cYYPJPSSFFPFKKXYrz�����������������������������������������������������������������������������ƽ���������������ý�������������������������������������������ynga\v���������������naaYO=4,%%,3<DOTBOOB<<6993),/66<<DTa�����vnannnbnn��������yy������������������yyv�zpp^E<<<EW\pvzpvv�zzrmw����������zrnga\aaaaYYOHHF;JHEFM;;;PYrz����ø������������������������������������������������������������������������н��������ƽ����ƽ����������ó�������������������¼���������zpgaa[gz�����ų���������vnaYTA6*,,6DOWWOODB6666/))%.6<EOELav�����vnnvvvnnv��������vz�����nvnvvyv�������vnnnnnnnv�vnOOLLOanwz�z�z��yznnw��������wznrnnag\YPPPOEE=;FEHPMF;;Xcmz�����Ƹ�����������������������������������������������������������������������������������̽������ƽ������ó���������������������¼������zmaang\ny�������®���������ynYE<4)37>TbbWOE64.3)).)),4EDEDbnvnv�����������������vnvvzy���nbWWbnnnv���vvnaaaanWTavnanpnnngpppw��������mn������zzrwnamvng\YPEEHPPHEF?=?VPFFFXZs��������ð����������������������������������������������������������������������������������ƽ������������Ѽ�����������������������̼�����rYRab[an��������ż����������vnWOD9%*4=OWabaO<,%%%,-.,4<BEOWbnvbn�������������zvvnvvnnpynWWDEOObaanvvnnabWOYYOOLTaaYanrz��������������zwz����zwrnaaanraSSHE=EHPYPEHFEFP\ZYYZZs�������н���{��������������������������������������������������������������������Ľ������������������������Ƽ�������ƽ��Ƽ�����������Ź��wgYW\Wanz��������ϻ������������nbOD</.<EaaabnOE./4<<BDDWannnanv������������vnnababaWb]]WTOO<D<EOTWannnnagWREEOET^aWT^nv�����������������������nnaaacrmcOEH==HYYaYPPJPYS\\\lmcs{������İ������������������������������������������������������������������������ƽ������������������������ƽ������������ѽ����������ѹ��papgbgnv���������ȼ�������������nWWEBLWbavnpnaO6).BEOLOWWapvanp������������pn]]]Wbb]TDDEB<<<<<9DOWbnnnnaWWOELAOYTYOY^av����y�����������������raaa\\ca\\YPPPEPYmacaa\YYSY\\aluos������é��������������������������������������������������������������������������ѽ������������������������ý�����������ƽ���������Ѽ��mnzyvvzz����������·������������vkWOObnvvv�vWOD6%/DOWWWabbnvanp�������������vnWTOTWWbTB6666666B<BHWnnnanaWOOYLLWWOOOTanz���������������������wnYY\\YYWORPS\YYahzwwmgahc\YP\\cmms�����������������������������������������������������������������������������������ƽ����������������������������������������¯������Ũ�yp��y�������������������Ź������vnnanv�����bOD<)%36<EOWb]nakbvvvany�������������p]OLBBDWTL</.)466BEEOOOWWbWTbOWO\OOOYOOOWanz���wpz���������������zna\ROOOOORSagrww��zwrwmrmmYYYYgacw���������������������������������������������������������������������������������������ƽ������������������������������������¼������ڼ����z���������������������˼���������vy������vWOO9./6<EEDWabknnabannWny������������vn]D9963<BB6%39<BD<<DOOOOILOOOWYWOYYOAELYarr��wnny���������������vpgWOOEEOY\awz����zzzwrrrwnaYag\amx����������������ƽ����������������������������������������������������������������������������������������������������������̹�������Ƽ����������������������������������������������aWWLOEEOWWbjnnnvvnWbakan����������vnnT<6,,%.44.%/6<A<96>ODDDDB<IWbY\OOTOE<<OYkp��wagwz��������������wwgWH==<OY\g���������wmrrrwhaaa\\ccw��������������ƽ�������������������������������������������Ľ���������������������������������������������������������������ż�������ż�����������zzyy������������������������������nvnaaOWWnvppvv��nnnnbavy�������yvnnnnaWI9,)%,%%)./66666<6<BBDDOOWbROa^O=6=EPkrvwn\nzvz��������������pn\aHE<HOYh����������rrrrraaa\Y\S\cZmmx{��������ƽ����������������ƽ��������������������ĵƸ�ƽ�������������������������������������������������������������������¼�������¼�������wwnav�������������������¨�������������vaavy�y��ynnnanvy�����vnaWWWWW]O<.),)%%)644,)))6<DIIOORORYnnO=EOOEYkananz��z��������������zggn\RO?Paw����������zwzrrnnghZS\g\SZlms�������ƽ�����������������������������������������������������������������������������������������������������������������ż���������¼�����pkaapnnnv�����������������ż������������������������vanvy���vkbOOOWW]TB9/)%%%,,%))4<DDOIOOI\annaOW^aaannanw������������������wnmngaRW\nz�������������wrrnrm\Yac\\\Zmw�����Ƹƽ�����������������������������������������������������������������������������������������������������������������Ѽ�����������ż���nWWabbanv��������������ż�ż����������Ů������y�������vWnnyynvvnnb]OOWWbWTL6/),%,/,6<<EDO[agaaaanvvwpz�������������������zz�wmnng\agr�������������z��zzmah\amh\\hr�������ƽ��Ʃ���������������������������������������ĵ�����������������������������������������������������������������������������������ų��kWWWWTap���������������˼��������������®�����������nOabnnnnvvnvnnaOObbbWWO</,%%%,6<DIRaW]nwwpy��������������z�������yzwzrmnranwzz�����������������zzmmrwzhchrz����������ļ����������������������������������������ĵ�����������������������������������������������������������������������������������³��nbROW^av����������������˼�������������˼����������vbWaW]babbnnnbkbabnnkaWO<6)%6BDROOYnv�����������������������yvwwzzzwww�����������������������zz�zwzmr�z����������������������������������������������������İ���������������������������������������������������������������������������������ż����pnbWkanv����������������żŹ�����������ϼ�������yyvvvvabWOEDLWOWnnbb]bannnnnbWO</-

.9AELOTnv���������¼�����������zzpgrw��������������������������������zzzzz�������������������������������������������������������������������������������������������������������������������������������ų������¼�����vpnnpnv�����������������ϼ�ű������������±����vnnnnvnbOE<69DOWaaaWWanvnnnynWOWL6/,,,


)6EELOWn�������������¹���������zzngmn������������������������������������z��������������İ���������������������������������������������������������������������������������������������������������������Ŵ�����ż��������zyy����������������������˹�������������ż���vnaWObnnWO<64.<EOWWabbnnvn�nnWaWO<66.)



%//DO[Wgv�������������¹���������zza^Yg��������¼�������������Ƽ������������������������������������������������������������������ý�ļ����Ƹ���������������������������������������������������������������Ƽ�����ż��������������������������������ű��������������Ϸ�nWWETWaWOO6,4/49DDOannnnvvyyvnbaaaO<664)).))/6DObba������������ż�³�������zvYWYn��������̼�������������ƽ�ó��������������������������Ľ�����������������������������������Ƹƽ������Ѹ���ƽ����������������������������������������������������������̳����ż���������������������������������ż�������������ϱ�vbOOEDDOE<O/,.),9DDOWnnvvvvvpyvvvannnO<6466,
%./6,),.9DOabbnv�����������ż����������vpna\Yn��������̼��������������������ü��������������������������Ľ����������������������������������ý����������ƽ����������������������������������������������������������Ƽ������¹�����������ų�������������������³������������¨�nWTE6699D6D,-%)-4<DOWnnnnnnnnyvvypvnnO9966,%,/,,4.,6BObWabg�����������ű����������vvnnbaw���������®������������������������������������������������������������������������������������������������Ƴ�����������������������������������������������������������������ų�������������������������������ϼ����������������vbTD4/))6DE,,4BWb]aavvnvy��vvaOB<6.,..366666<<DEOObankn������������������������zwprz����������®�����ó�����������������������������������������������������������������������������������������ó�����������������������������������������������������������������³���������������������������������ű��������������vbO96%%<O))4<OWbWWnnnn����������v]O<<9<<<DD<96<OOTT]anvnvv���������������������������z������������¯�����½�����������������������������������������������������������������������������������������ƹ��������ü������������������������������������������������������������������������������������������¹�ż��������ű�nWB6)%6O)<LOWaWaaanv�����������pWELODOOLOO=<EObnnnv�����������������������������������������Ƽ���Ƹ��Ƽ��������������������������������������������������������������������������������������������������Ƴ�������������������������������������������������������������������������������������������˼��ż������˱��nOB6)/9/.-4<LTWaYWOav�y�����baOWWaabbaWOOavz������������������nnny�������������������������������¼����������������������������������������������������������������������������������������������������Ƽ���������������������������������������������������������������������������������������������ż��¼��˱��vaO<<)%/994%%%/9BBOOOOOnvvy�����vnabavnvnvbbbbn�������������������nnny������������������������̼���������������������������������������������������������������������������������������������������������½����������������������������������������������������������������������������������������������ż����������nnWWD6.%BB4,%.4946=<OWavvnvvy����yvvvvv�v��vnnv������������¹�����vav�������������������������¼��������������������������������������������������������������������������������������������������������ü����������������������������������������������������������������������������������������������¼����������vnaaWO</)%DE9,),..46DWObannny���������������v���������������¤����v��������������������������Ѽ�������������������������������������������������������������������������������������������������������Ƽ��������������������������������������������������������������������������������������������Ź�����������vnbWOOE9,%,)%%%<</.%-66<DWabnnpvvvvnp��������������������¼��������ű����������������������������������������������������������������������������������������������������������������������������������������ƽ���Ƴ���������������������������������������������������������������������������������������ϼ������������nanWWOOB6,.64,%,%9.4%%%)4<EOWaabnvvvvnnp��������������¹��������������ų����������������������������������������������������������������������������������������������������������������������������������������ѽ��������������������������������������������������������������������������������������������ű����������znaaOODOO<<6<<99/%%4/)%%%49BTOOWabnnnnnp�����������������������������ϼ������������������������������������������������������������������������������������������������������������������������������������������Ƴ��������¹���������������������������������������������������������������������������������³�����yvabOO<<6EOEOOEDOT9),44.,,<DLDTTTaan]bn����������������������������ż���±�����¼�ż�������������������������������������������������������������������������������������������������������ƽ������������������ư��������ƹ������Ƴ�����������������������������������������������������������������������˼�¨���nbaaaWWDEE666EWaaabbWbE/%46)%6<BDOOOWabbaWn����������������������������³���¼������������������������������������������������������������������������������������������������������������������ƽ����������������ѽ���������ƺ����������������������������������������������������������������������������������ű���vaOOLOE<66/<<WbnnanannT46.
66<<BLODOWWWWav���������������������������¹���������������������������¼�����������������������������������������������Ƽ�����������������������������������������ü�����������������ƹ��������̼������������������������Ƽ������������������������������������������������������żŮ��v]LDOBEE</46EWbnvvnvvnaTBD/.,9<D<EET]Wbny������������������������ż����������������������������ѹ�´����������������������������������������������ù���������������������������������������ƺ�Ƽ����������������ï���������̽�������������������ż�����������������������������������������������������������ϼ���vYDLDOEE<69BOanv�vnWTTb
%%,9<<<ETTbav�����������������������ż�������ż���������������������ż�������������������������������������������������ó������������������������������������ѽ�����ü�������������ƽ����������Ƽ�����zz�����������ų������������������������������������������������������������ϼ���vaTTOEEOOEEOObnv����nWOOan%%%).4/9BLWanv�������������������ϼ�����������˼������������������������ż��������������������������������������Ƴ��������������������������������������������ƽ��������ý����������ó�����������������zzz���������ų�������������������������������������������������������������ż���nbYTEEOOOOWWbnv����aWWOOW,%%-%%/69BEOanvv��������������������ż�������������������������ż�������������������������������������������������é��������������������������������������������Ѽô������ü����ƹ��������������������������������������������������������������������������������������������������±����vpnbWWbbbWabn����nbaOOT3/
%,.),,,66<OWnnn�������������������ż������������Ź����������ϼ�������������������������������������������������ڹ�����������������������������������������������ý������Ƽ������������������������������������������������������������������������������������������������������ϼ���������ynnnvnnnnnn����vnbWWO<6%%--4/../-9<LOaanv��������������������������������Ź������żż���������������������������������������������������ѹ������������������������������������������������ƽ������ý����������������������������������������������������������������������������������������������������ż���¨���������vn����vnWbWD4,%%),.6/.%))))44,-.)49OEOWav����v���������������������������ϼ�ż¼�������������������������������������������������������ѽ����������������������������������������������������ýƼ³�������������������������������������������������������������������������������������������������ű�����ż¹����������������vnnWWOD%)4<BTE<4,-,)%))-,4.,4<<WanvpnaWanv��vnn������������������ż�����������¹����������������������������������������������ƽ����������������������������������������������������Ѽ����������������������������������ż����������������������������¼����������������������������������ϱ������ż��������Ż��������vvbWO<%,6<OWOA6.,%).464,6<OWnnnvnbWOWWWannnbWbv����������������ϼ����������ż�����������������������������������������������¼�����������������������������������������������������ú�����������������������zrrz�������³���w�y�����������������ż���������������������������������ż���ż�����������������˻��������vnvvnbE6%,46DOOE44/%/64.,.9OWWnnnnbWOWOEOWWWOOOavzvv������������ż����������±���������������������������������������������¹���������������������������������ƽ�����Ƽ������������ƹ�����������������������zrwz������Ѽ���zngn����������������Ź��������������ż����������������Ź�����ż������������������·������vnv��nWE%.4<B<64,,.,)%.6<DObWaaabOEDDB<D<D<BOWnvnvv������������¼���������¼�������������������������������������������ƽ����������������������������������Ƽ���������������������ó�Ƴ��������������������zw��������ų���nnnny��������������ϳ�����������ϼ������������������ż���������������������������»������yvv�����nb),,)%%%%%%%,4<DOOWWnbODEDD<<<<<DDTWaWan���������������ϼ���¼���ű������������������������������������̼���ѳ����������������������������������Ƽ�������������������������Ѽ������������������������������Ƽ���pvpv����������������ϼ���������˹�����������������ż�����������������������������ŷ���������������y
%-6DOOOWbWWODOO<D<6669BLLEOnnvv���������������������ż������������������������������������ż�¼��������Ƽ������������������������ƽ����������������������������ƹ�������������ѽ�������������������zzpvz����������������·�������˼���������������ż����¹�������������������������˷�����������������%)-6DEOWWWWabOWD<<<66/.66636OWavn���������������������ż�����������������������������������¼������������������������������������ù������zzzzz������������������ƽ���������������¹������������������wppy����������������»���ż��¼�������������ϼ���ż���������������������������ռ������������������

),6<DODOOEWWaabE<D</))..,.46EWan�����������������������ż��������������������������������Ѽ������������������������������������ù�������zzrwwz�����������������Ƽ����������������ڽ�����������������vvpnp���������������ż¼���¼�������������������������������������������������ű������������������
%46IED<DEOObnaWODB6)%))44/<Wn����������������������������������������������¼���������ڼƼ���������������������������������½�����zz�z�zzwpz������������������Ƽ�����������������Ѽ����������������ypnvz�����������������ż�¼�����������vv����������������������������������������������������������
)).4BB<9BEWbannaO9.-//%334Dan�������������������������������������������Ź���������¼�ż��������������������������������ڼ����zznrzv�zwvpz�������������������Ѽ�����¹�������������Ƴ���������������wvy�����������������ټ�������������vnnnvv����������������������������������ϻ�������������������


%,44<9<9BOannnbWE6-)/94%%6<EWnn������������������������������������������Ź����������������������������������w�����������Ѽ�����wrnz���wrnz�������������������˼��������������������Ѽ������������������������������������ϼ������������nnvvvv������������������������������������»��������������

%-/46646<OaaaWODB4%)9E9%%))/6OOObv�����������������������ϼ��������������¼������������������������������������rnrr���������Ѽ������rwz�����ww���������������������Ѽ���������������������Ũ�����������������������������������ˮ������������pvyy��v���������������������������������������ϻ������������
%%%,449/46DIEEE<444-.4<<44/9DOWWWav�������������������ż¼�����ż����ż����������������������������������������znaaYgn������Ѽ����zzw����������������������������������ż��¼���������������Ƴ������������ż��������������������ϼ�����������������������������������������������������������������������%,,%).4/-./46449<,%%),-449EEEOnbWObnv�����������������ż���������������������������������������������������������zm\OERaw���������wwzrrz���������������������������ż����ż��������������������̼������¼�������Ź�����������������Ѽ�����������������������������������������������������������������������%%,,4.39664/.))43-%%,),-/))%%%%)4=EEObnvnvvy����������������������������������������������������������z�����������������w^HHPan��������pgmwwn���������Ƽ�����������������ż����������������������������ż��������������ŷ�����������������¨����������������������������������������������������������������������),..DDELLLB9/,,%)-%%%,%)%%,6DWObn��������������nnnnv���������������������������������������������zz���������������wzpYHEYYaw������m\O\nwr�����������������������������ż�����������������������������Ź������������±�����������������Ů������·��żű��������������������������������������������������������-3<BOabaWTL964./,-4/%%
)--,<EWbanv�������������nWOObabnnnnvvvvav������������������������������������w���vvz��������yngaYRSRYamw���znWOORarr�����������������������������������������������������������Ź������������¼�����������������ϼ�������������ϼ���������������������������������������������������ŷ���,6BLLWnnnba]D<966666/),%)%%
%/66OWnnv������������vnWOIWWWaWaWnbbbWbnvv���������������������������������w��vnpz��������vngYaYYY\amz���naWER\pzw���������������������������Ѽ�����������������������������ż������������˷������������������ų�������������ż��������������������������������������������������±����%%/<DTOannnnnaTEB66<<<4/64/.),%-6EDWWnv�������������vabOOITTTOOOOWWWOOWabn����������z���������������������zz�papv��������va\Ygga\aap��z�raWORaw������������Ƽ�������Ѽ�����Ƽ��������Ѽ��̼���������������ż�������������¨������������������³�������������ż�����������ż�¹�����Ż���������������������������������%%4AOWWnvnnnnnTODB<OEO<<<64)%3.,%%4<OOWWny�������������vaWWEDLOLO<<DOTOOOOWWav�yvvvy���zvn���������������zywnvwnagp�z������pa[aagaaaanv�vygYWEYgwzw���������¼��������®����ż���������¼¼����������������ż����¼�������·���������������ϼ�����������������������������ű�����������������������������������˱���y���),6LWkknvnnnnbOTLLOWYbOED<94,.63-%./<EWWWWnvz�����������nabWOIOOLO<6<EOTOEOWWavvnananv�zvn��y����z����zvnanpa\bnvv�����ypaaaa[gnnagpvpvaYOEY\npm������������������³����������������³�����������������ѹ���������Ż¼������zv���������±��������������������������ż��������������������������������������±����y��),<O]kbnvvnnnaILLOWnnnaOODB9.6B9//,,%6<OWWWaannpvv����������nbannbOOOOL96<OTTWOWbWavd[YgWYn�vvyvvppyyzzrz���zvnanpbRRgppv����vpanngnvpra\annn\YWRYYggnvz����������������������������������������������������Ƽ��������������������vnv����¼��������������������������������������������������������Ż�����������������vv