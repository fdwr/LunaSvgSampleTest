��  ����������˼����˼�����ڼ��ڼ��ڼ�����`$-9-999B9B9BBBPBPBPPPBPBBBBBBBBBBBBBBNBNBNNN\N\N\\\\\\\\ffffffffffffftftfttjtjtjtj�t�������������tttttttttttttt~�����������������~�~�~�~Zf�@@t�������������������hZ~�������������ڵ����������������������S���������z��S�����mttttttttttjtjtjjj\j\jf\f\\\\\\\\\\\\\!!!8���������������������������˼��ڼ��w��`(-03UK<<<G<GB;B;B6B;;;B;BBBBBGBGBGGGGGGNGNGNNNNNUNUU\UaUaafffqmqqqmqmggjgjcjjjjjnjwn|t|����w�||ttttttxtxtxxxxxxx���������������~�~~~~~~~==8�D~�~z=8@81X~��������X=�~�~�~�~�������̘��������������������q����������M�X�������tnnnnjnjnjjjjjcjcjcccccccc\c\\\\\U\UUi���������������ü����������ڼ���ڼ�����`-333aNa7<B<;B;;;B6B;;;;;B;B;BBBBBGBGGGGNGNGNNNUNUNUUUUZUaZfZfmfmmqfgfggngjcjjjjjnjwnww|||�|w|w|n|ntttttttxtxtxtx�����������������~~~~~~~~~z#�#8@1=�~�~�X=d�������QD��~�~�~��������Ҙ�������������������q����������Hw�B�������mnnnnnjnjnjnjjjcjcjccccacaNG\\U\U\UUU!!q���������������ü�����������Ҽ���ڼ�����`-339_�e<C<7<;76;666;6;;B;B;BBBBBGBGGGGGGGGNGNNNNNUNUNUUaZfafmfmmqfqmggcgccccjcjjjnntn|x|x|w�w|ntntttttttxtxtxxxxx���������������~~~~~~~~~��1�JZt~~~~~~~~~7k������Qq�~~~~~~~������ּ�������������������q�����������+��S��������jnjnjnjjjjjcjcccccccccc\c\NG\\U\U\UUp7q���������������ü�������Ҽ���ü���ڼ�����`(3939<97<77;7};666;6;;;;;;B;BBBBBBBGBGGGGNGNNNNNUNUNZUZZZZfafgmmfafgagaccccjcjjjnnwn|t|x|wwwwnwntntntttttttttxtx|����������������~~~~~~~~�x@�Jf~~~~~~~~~�z*k�����`X��~~~~~~�����ּû�����������������q�����������w�`���������mnnjnjnjjjjjcjcccccc\c\ca\\'UU\U\UUNq�����������������������������Ҽ����ڼ�����`(999C97<77076Y6066666;6;;B;BBBBBBBGBGGGGGGGGNGNNNNNUNZUaZfgfgmmfmfgacgccccccccjcjnntttx|t|nwjnntntntttttttttxtx|����������������~x~x~x~~~~~J�Zt~~~~~~~~~~�Dst�����8�~~~~~~~~������˻����������������q�����������H+��`����������njjjjjjncj�ȩ��ccccc\c\c\\<5\U\UUNUq����������������ü�������Ҽ���ü����Ἴ����`..9393373776060666;6;6;;;;;;B;BBBBBBBGBGGGGNGNNNNNZNZUZZaaagfgfZfaaaac\c\ccccjgjnntn|x|n|nwwwnnnnntntntntttttt|||��������������~x~x~x~��~~~{�Qx~~~~~~~~~���XX�����Dx�~~~~~~~�������ҥ��������������q������������J��m����������mnjnjjjjjc�*o7u�c\c\c\\\UaN2UUUUUUNJ�����������������ü�����������ڼ�����Ἴ�����!93933030000006066666;6;6;;B;BBBBBBBGBGGGGGGGGNGNNNUUaUacagmgfafaa\ac\c\cccccccgnmtmxtxtnwjwjnjnntntntntttttttt|��������������xxxxxx~�@N�xxp�M~~~~~~~~~~~��D�D�����D~~~~~~~x~x�����ҥ��������������[�����������xBǬ�J���������vjjjcjcjc�2*}cc\c\c\\\U\!\UUUUNU4��������������������������ڼ���˼�����弼�����.3.333-30-006066666;6;6;;;;;;B;B9BBBBBGBGGGGNGNNNUUZUa\agagaZfZaZa\\\\c\c\cccgngnmttntnwnwjnnnnnnnnnntntntntt||�|����������|��xx~x~x~��x~X��=~~~~~~~~~~���|aQ�����k#X~~~~~~x~x����֥�������������J������������7���X����������njjjcjcj]>-B7-Pc\\\\\U\U\U.UUUUNUN4����������ü������ü����ݠ�Ҽ���˼�����弼�����/3(3----0-00000�6066666;6;;;;B;BB3VBBGBGGGGGGGGNNN\U\\acgcaafZaUa\\\\c\c\cccgcmgmxmxmnnjnjjjnjnjnjnntntntnt�tt||�������������xxxxxxxxxxxx8��@~x~xX*@1d~~���Dh������d@8DXt~x~xx�����ƞ�����������q�������������`���`���������mcjcjcccp�V\\j�\c\\\\\U\U\!UUUNUNU�������������������ü����F��˼��ڼ������Ἴ�����Y(3(3----0-0-0T2T66666;6;;;;;;;;B;!)VIBGBGBGGGGNNUUU\\acacaZaZZZaU\U\\\\\c\cagggmtmtmnnnnjnjnjnjnnnnnnnnnntn|n|w������������|xtxtxxxxxx~xqeږXx~x=R~~~X=����L�Q����~xdLtoX8Xx~x�����ƞ�����������+�������������(-����XBS������vjcjcjccc����т\\\\U\U\UUJ'UZUUNUNq����������ü�������ü���h�ڼ���ڼ������Ἴü���p$(-----}Y0-00�u�06066666;6;;;;B;B(IGBGBGGGGGNGNUV\\ccca\aUZUaU\U\\\\\c\c\cggmmmqmgmngjjjjjjjjjnjnjnnnntntntn������������|xtxxxxxxxxxxx=��<xxx7x~x~x~mJ���hkL�����~xXD|���=_x����ֻ�����������Jh�������������z0ZZPu��ǹ�Xq�����dcccccccc���\c\g\\\U\U\U*JUNUNNNNJ����������ü��������ü��V�ڼ���Ҽ������ڼ��ü���((-(-----0->0�060666;6;6;;;;;;B;$R;V\BGBGNNNUVU\c\caUaUZZZUUU\U\U\\\\acagfgfqmggngjnjjjjjnjnjnjnnnnnnnnnn|w�|�������||||ttxtxtxt�txmeڸ@xxXR~x~x~x~�Q���D=����~x=_~R���ȁ=���Ǽ�����������q�������������کU660(IǬ����q����mcccU8c\c\c\\\\\U\U\UUU'GUUUNZNUN+�����ü��������������ü�!��Ҽ���˼������Ҽ��˼���/(-(-----0->f0000606066666;6;;B;((-P_NNGNNVVVc]c\\\UZNZNUU\U\U\\\\\cagfmmqmgmggccjcjcjjjjjjjnjnjnjnnnn|w�|�������|�||ttxtxtxtxxxxM��emxx#gxxxxxxxx�DY�b2�����Dmxxx_���Ȼ_���û�������������������������Y0!+�����X�����ccUX8cc\c\c\\\\\U\U\G'JUNUNNNNNGq����������ü����������ó$�������˼������˼��˼���p!(((-(-----0-006060666;6;6;;;;;;B;3*-?mINVNVcVc\U\UZUZNUUUUUU\U\U\\aaaafmfgaggcgjcjcjjjjjjjnjnjnjn�ȩ��ww|������w�w|t|ttttttttxtX�کRtxR.nxxxxxxx���`@g*��z_8xxxxtxZ�������˻���������4h����������������X�����J����cUQ�\c\c\\g\\U\U\UU'<UUUUNUNUNUNJ�����ü���������������å!!V�ڼ����˼������˼���˼���((-(-----0-0000006066666;6;6;;B;B;B7#0zVVV]V]V\VUUNUNUNUNUU\U\U\\a\fafqfmfggccccccjcjcjjjjjjjjjnj�*o7u�|��������w|ttttttttttxtd���Itxx8aaxxxxxxxx����a*=88Z�xxxxxxx_���Υp��å�������io����������������ǚ����J����W�.c\c\c\\\\\U\U@GUUNUNNNNNGNG������ü�������������Ҽ�!!!w�������μ�����弼���˼���J(((-(-(-----0-006066666;6;6;;;;;;B;BB3-lPVV]VUVUUUUNUNUNUUUUUU\UaZaafffafgagaccccjcjcjjjjjjjnjnj�2*}w|������w|w|ntnttttttttN��ZtxtxQ�Dxtxtxtx|�����L8}�|xtxtxtxtxZ�������å�������z�����������������ǚ����J��qg�\\\a\\\U\U\U8a'UUUUNUNUNNNGNJ���������������������ˑ!!!�ڼ�����μ�����弼���˼�˒�(-(-(-----0-0000006066666;6;6;;B;BBBB7#!xV]VNVNNNNNNNNNUNUNUU\U\Uaafffmfgacaccccccccccjcjcjjjjjj]>-B7-P|x�x���|�w|ntnttttttttI��Ztxtxcw�Dtxtxtxxx������*�|xtxtxtxtxtx7�����ݸ�������4������������������ǚZX���J�q*��@c\\\\\\gU\UL�QCUNUNNNGNGNGGG������������ü��������X!!!��������������鼼���Ҽ�ˣ�J((((-(-----0-0-006066666;6;6;;;;;;B;IBI:.w]PNNNNNNNNNNNUNUNUUUUZUaZfZfZfaaaac\c\c\ccccjcjcjjjjjjj|�V\\j�t|���|w|wwnwntntntntnR��Zttttt@��Dttttttx|������LT�|tttttttttttR����ˬ������iU�������������������ǚa���w`**2�hD\\\U\U\U\U8àGUNUNUNUNNNGNGNJ������������ü�������{!!!!!��������������弼���ڼ�����((-(---�-0-0-0000006066666;6;;;;B;BBIIPIPV;j]NVNNGGGGNGNNNNNNNUNUUaZfafgfaa\ac\c\ccccccccccccjcjcjjj����ѓ|x�x�x|nwnwntntntntn_��Dtttttt<�ictttttxtx|�����w*ZxtttttttttttM���˼�������!$0��������������������ǃZX���2%w�hD\\\\U\U\U@ww?UNUNNNGNGNGGGGG�������������ü�����ݐ!!!!��������������Ἴ����μ�ˣ�p!((6(-P2T---0-00006066666;6;;;;;;;;IBIIPPPVPNINIGNGGNGNNNNNUNUNUUZZZZaafZaZa\\\\\\c\c\c\ccccj��cjjjjj���n|t|x�x|wwwwnnnnnnnnn_��Mtn�wtnci�<tttttttt||||����?sZttttntntntntD��ì�����47:0(����������������������+77�����hN\U\U\UUUU.GUNUNUNNNNNGNGGGGJ�������������ü�����!!!$!!�������ڼ������Ҽ�����μ��Ғ�/$:f-(�u�--0-000000006066666;6;;;;I;PIPPPVPNPNIGGGGGGGGfTNNNNNNNZNaUagfZfZa\\\\\\c\c\cccccccj?Ljcjcjcjnntttxxxtx|nwjnjnjnjnngJXZtnt|tnt8ǖRttttttttt||�����pX�Zttttntntntn=���ˬ����477C0$!o���������������������`a��`@@��hN\\U\U\UU#<NUNUNNNGNGNGGGGGGG��������������ü�����7�P!!!!$!!���������������˼�����ڼ��ҵ�p!(((((�(-----0-00006066666;6;;;;BBBBPIPVPIIIIGIGBGGGGNK:\|tpfZZUZUaaaZZZaUaU\U\\\\\c\c\c\ccp��pjcjcjnnnntxxx|t|nwnwjnnnnnnn*@cnnnnnntce�<ntntnt��ntn|w���w|?��Zntntntntnn[{��ˬ���i7;6H(!��������������������ǤZw�`*%g�o<\U\UUUU*GUUNUNUNNNGNGNGGGGBGB�������������������!!!!$$$!�������������弼�����弼��Ғ�/($((-(-----0-000000606066666�6B;BBPIPVPIPIIGBGBGGGGGG*H_aUa\aUaZaU\U\U\\\\\c\c\c\cccc��ccccjcjgnmxtxxxtnnjnjjjnjnjZMjnjnnnntn8ǖNtntnt|@N|n|w�����wpX��Zntntntntn���һ����x(0$o���������������������Z`�`**U�hDU\U\UU9'NUNNNNNGNGNGGGGGGGGGi�������������ü˘�7!!$!$!!������ڼ������ڼ�������μ��ҵ�v!((((-(-(-----0-006060666;6!0jP\ZcBIIPBIIIBIBBGBGBGGGC�UaUZZZUZU\U\U\U\\\\\\\c\c\c\ccccjcjgnmttxxxtnnnnjnjnjnj2@ZjnnnnnnnnZ��Innnnnnn��nnn|w��|www7��7nnnnnnnn�����ì��Pv-!���������������������BhJ�J**%al5\UUUU8*JUNUNU'JJZZMM!1<GBGBG��������������üX!!!!$%$!!!��������������ü�������ڼ���Ғ�/$((-(-(-----0-000000606066%-$->boBPIIBBBBGBGBGGG?.7*!n\aUZNUU\U\U\U\\\\\\\c\c\cccccccccccmnmxqxmxtnnjjjjjjjZ{UjjjnjnjnjnF�Znjnjnjnnnnnn|w����|wwM���Gnjnjnj������ì��Z~>��������������������Ja`�``B8�8U\UG;�'UNNN?;�������Ҹe'GBGB+�������������Ҽ>!!!!!!$!!!!�����ڼ������ڼ������������ҵ�v!(((((-(-------0-00606066!0bbI;IBBBBBBGBGBGGGGN9*maUZUZUUUUUUU\U\U\U\\\\\\\c\c\c\cc�pnmtmxmxtnnnnjjjjj^�Njnjnjnjnjn2�Snnnnnnnnnnnnnnww|�|wwww=��7nnnnjn�����ݻ��diz��������������������JZm�S���J.1UJ't�LJNUNGw������������WGBBJ��������������s!!$!!!!!!�������������ü���������ü���ڒ�/($((-()!MMQZZSS7!)-0060%)0737bBBBBBBBGBGBGGGGGGGN<2828\UUNUNUNUNUU\U\U\U\\\\\\\c\c\cccccgcmmmqqxmnmngjjjjjS�<jjjjjjjjjjU�Sjjnjnjnjnjnnnjwn|t|x|nwj2���Gjnjnj�����ô�v�>7�%*�������������������BZ`�J����qG'Q���'NNN?|��tJ!!!%!8����*BBp������������Ҭ!!!!!!!!!e���μ������ڼ����������μ���ڣ�Y$(((Q����������ܚo%60676;;B3%\;B;B;BBBBBGBGBGGGNUNUVU\UUUZNUNUNUUUUUUUU\U\U\\\\\\\\\c\cacagmmmxmngngjjjjjG��Gjjjjjjjjj]JSnjnjnjnjnjnjnjnjwn|x|nwnw@���8njnj2���˼���T�Z������������������hw�B�����k����DNUN?o��?5BNGGGGB.���]B;��������������{!V;!!!!!!��ּ�������ü����������Ҽ����ǘ�$X����������������t%067;<;BGB;I;B;;;B;B;BBBBBhBGBGGGGGNNVVVUNNNNNNNNUNUNUUUU\U\U\\\\\\\\\c\c\cggmmmqqqmggccjcjYt�Fjjjjjjjjjj*2jjjjjjjjjjjjjjjjjjtttxtnnjPh��7jjj^�����ü�v���>**m�����������������77+��B���������DNNNG.�|!GGGGGGGGGB'��g;BB��������������w!!?5!!!���������ڼ�����������Ҽ����ڃ�J3������iM!!!Fcl�����Q7;7;BBI;B;B;B;;;;;B;B;BBV}BBBGBGNNVNVUNUNNNNNNUNUNU\UUUUUU\U\U\U\\\\\\\\agagfqfqmggggjcjc2��8jjjjjjjjj*Gjjjjj�jjjjjjjjjnjjnntxtnnnnPh��Jjj^�����˼��T���o*%8�����������������hwǬB�������|=NUNN5o|9NGGGGTGBGBG3�]B;S��������������{!!!.a!!!!M�������弼�����������Ҽ�����i�T���a3$((-------)o���Q<;<G<;B;;6;6;;;;B;B;BBB<!YUBcuNNVNVNVNNNGNGNNNNNNN<QgtuZ\U\U\U\\�p\\\\\cagfqqqmgmggcccc]o�zVcjcjcjjj22jjjjja2ajjj�wjjjjjjjtttxtnnj\h��Zj2�������˴vT����*?g�����������������Z+Ǭwi������c5NNNGN!g9GGGGGGGGGBGB;�!;B���������������3!!.!!�������Ҽ������������Ҽ�����VT��X!$((((((-(-----0()B��N<B<;;;B6B6;;;;;;;;B;B;.$-(Kc\PNNNNNNNGNNNNNUNU!-;cuUUUU\U\U\U\\\\aafffqfgfgac\cccG��FcjcjcjjjUDGjjjjj�u�jjjwjjjjjjjnntxtnnnn\h��J]t�������ˎ�J���hJE�����������������aX��B�������ZNNttNG@!NGGGGGGBGBGB;Q�Q;B;��������ü�����!!!!!!������ڼ�������������Ҽ�����]��$$($($((-(-----0-030.e�'<;<;766666;6;6;;B;B;B%!!$:ccNNGGGGNGNGNNNN'!!$(�hU\U\U\U\\\\\\fffqmqfgacccccc8��1ccccjcjYXQccjjjjj�jjjjjjjjjjjjjtttxtnnjPh��78��������B�B��ȗh�����������������h�ǍJ�������NNU?LN<<GGGGGTG*!7QJ!;B;;��������ü����?!7������ü�������������Ҽ����`�Ti$($($((((((-(----3737.SS07;76;6;6;6;6;;;;;;B;B;BB;$BVGNGGNGNGNNNNNNNUN<-gnUUUUU\U\U\Uaafffmfaagac\c\c8�@cccjcjcD�*cjjjjjjjjjjjjjjjjjjjnntttnnnnPh��8<������饨�B����7u�����������������VZX�`��������^Nh��a1GGGGBGBGBB3***B;B;;;�������������Q!!h�����ּ��������������Ҽ���es4��/$$$$($($((-(----30379<<1!07606066666;6;6;;B;B;BBBBI:22225GGGGGGG\NGNGNGNNNNNN<818NUNUU\U\U\aaa�����nfgac\c\c]o�zNccccccG��@ccjcjcjcjcjcjjjjjjjjjtttxtnnj@��a<i�����>��������u����������������ڠZ�`��������^NNnnG!!GGGGGBGBGBBBBB;B;;;;������������Q{����ּ���������������Ҽ�û#�S��B$$$($($((((((-(3333979737606066666;6;6;;;;;;;;B;IIIIPIIBIGBGGGG6VRmuNNNNNNNUNUNUNUUUUUUUU�hj;%%-PP[a\a\\\\Qz�]c\c\ccc<�pIcjcjcjcjcjcjjjjjjjjjnntttnnnn@��32���ږ>t��������zh!5h������������������guAwi�������XUNNGG.GGBGBGBBMBBBB;B;;;;;���������üe�!!���ڼ����������������Ҽ��]e�S��J$$$$$$($($((-(3-339<9730!0000606066666;6;6;;;;B;IIPIPIIBIGBGGGG#<}aGNGNNNNNNNUNUNUNUU\81aa\a\\\\c@��!\cccccQi�pIccccccccccccjcjcjcjcjmtmxmngj1��2����]z����������ah>!66H$u�������������������EXB��������NGGGC@!GGGBGBGBBBBBBB;B;;6;���������üo{���ü����������������Ҽ��>��S��S$$$$$($($((((.(3.9393373!-00606066666;6;6;;;;;;BBIBPBIIIBBBBGB*!!'TaGNNNNNNNUNUNUNUUUU=@I==F`ZaZaU\U\\\8��*\\c\c\8��wI\ccccccccccjcjcjcjcjgnmtmngjg*�.|�Xh���uuuouhhZZZ7>�uuuu����������������ni�������UNGG<J!BGBGBBBBB;B;B;;;;;;6B���������æ?22!7��ü�����������������μ�X���Z��S$$$$$$$$($$!!+3933030000000006066666;6;6;;;;IB\BIBIBBBBGBGBGG96}GNGNNNNNNNNNUNUNUNZZagfafZaU\U\\\\8��8\c\c\c8��{Iccccc�pccccccccccccccmmmqmgg]%D���S!*8�����������������J%FhZ7E�uuohhaZZMBBM��7+X�������GNNG1|!GBGBGBBBBB;B;B;;;;6;J����������axu}��aJVQMa�������������˼�V���Z��B$$$$$$]g{������i8!(3--)-0-00006066666;6;6;;B;BBIBIBI;BBBBBBBGBGBG*.aGNN{{NNN\UUNhuaNZZaaaaaZZUaU\U\U\8ߚ@\\\\\VV��zU\c\c\c\c\c\cccccccccggmmmcN*J|����Z*\c\���ì��������������SB8��EJ������������igǗ7i������GNNI%�!BBBBBBB;B;BM;;;;;;;6i����������.�V�����ü�M����������弼�p���Z��B$$!o{������������ڸi<!0-0-00000000606666666;6B;IB�BI;BBBBBBBGBGBGGGB.***<GGGh@NcNN52\\PPP�c\\aca�nfcRgj;U\U1�{D\\\\\Jt��uNc\c\c\c\cccccccc]G8%]caS1.a�����L@Vc\c���ì�����������������iJB2�E���������������Jaaq�����NNNG!�3GBBBBBBB;B;B;;;;6;6;���������í4���whhhh���ÊS��������Ҽ�h����V��!B����������Ǽ�������Ҹe!-0-0-00006066666;6;6B;BBB�B;;;B;B;BBBBBBBGBGBGGGGGGNG��NNN*1Ua\aU=3GUUU\1�lJU\U\U@���uN\\\\\\\c\c\c\G1Fz��������˸�iM��wo%c\\\��ڬ����������������������J*�J�������������������������^INIJ�Q;BB;B;B;uu;;;;;;;6;6����������Xqi4J�����aJa�Ê`������μ�Q����S��>������������ô��hhhZZZJJJ)-000000006060666;6I;I;�;;;B;B;BBBBBBBGBGBGGGGGGGGGGGGNG91115NU\\\caUZNUNUUUU\U1�ZN\U\U\1���uN\\\\\\c\c\Y1F����������������ҊM*x8\c\\��ڬ������������������������J++�������������������������oNIIa�h7BBB;B;c@N\;;;6;6666B����������*#��������iM��p����鼼�J����S`t������������l.((((----!%!0-00006-%!ZZwwZZ!%;��B;;;;;B;B;BBBBBBBBBGBGBGGGGGGNGC!NNNNNUUUUa\aUZUZNUUUUUUU!�SUU\U\U!���uN\U\U\\\\Q*t��������������������ˊ*J\\\\��ά���������������������������iS�������������������������oPI5�æ*;B;B;;;��;;;;;6;6;6J���������wa.���������ÐM�p���Ἴ�V����S���å����ҥvSv��������lF!--((---!!000-?x�����Ƹ�����䩊\U;B;B;BBBBBBBBBGBGBGGGGGGGGGGNGNGNGNUU\c\UUNUNNNUNUNUN!�SUgU\U\h���h\U\U\\\\*t�����������������������˚<\\\\��ì������������������������������������������������������oVP!�ü%B;B;B;;;;6;6�666660i���������ih�����������Jt��Ҽ��a��ک��ҭ���ݻeV���������������h!!!!--)?������ǹ��������O-;;;;;;;;B;B;BBBBBBBGBGBGBGGGGNGNGNGNUU\U\UUUUNUNUNUNUNU�!UUUUUUh���hU\U\U\GM��������������������������Ñ?\U���ì������������������������������4�����������������������oPI]���M;;;;;;M;;;6;6;6;666����������VSQ�������������tJ�ü����ҩ��ß����Xe�������������������t!-----7�������Ǭ�����������-;6;;;;B;B;BBBBBBBGBGBGBGGt\GGGGaaGNVUVc\UUNNNNNNNNNNNS�1NUNUNNu���h\U\U\'�����������������������������Ñ?\��ᬬ�����������������������������JZ�����������������������oI%����ZB;;;;;;6;6;66606060����������S;��ü�ppww{����e���p���Iڵ����oX�����������������������t$--)������̨J3!Bi��������-;;;;;;;;B;B;BBBBBBBBBGBGUNGGGGaNaNNUV\\UUUUNNNNNNNUNDii<UNUNUBu���hUUUGM�������������������������������Á���Ƭ���������������������q��������gZ�����������������������oIe����S;;;;;;;;6;6;6666666�����������Xo�����ˠi]zښ���p�˖o�����L��������������������������F)�����J/-70<73-!J������?6;6;;;;B;B;BBBBBBBBBGBGBGGGGGGi�iNGVVVUVUNNGNNNNNNNN5�8NNNZNND���BUN'�������������������o@@JJ@@Q������è�ô����������������������`S������J�h�����������������������o!�����%;;;6;6;bO6660606060�������ðJt����������ڸeXs��p��I�����Z���������������������������鳧���i!)!0377)3?)60<����Ǘ-6;;;;;;;;;;B;B;BBBBBBBBBGBGBGGGGGNNVUNUNNGNNNNNNNNN*�*NNNUNU9{���%CW�����������������zSQ���������oI������ּ����������������������iB������g�a�����������������������o����ڼ;;;;6;6UB;6H6660606��������.J����������������eJ�p��o����Z���������������������������鳧���8)0-0!%73���B060<���Ǿ!66;6;6;;;;B;B;BBBBBBBBBGBGBGGGGGNNVVVNNGGNGNGNGNNNN8�5NNNNNN5���'h����������������tL��������������oD���üì���������������������J�Z�����J��Z�����������������������o����ڵ%B6;OO6666060606000S���˼��������������������ک.p�i����L���������������������������峗���h!---303<���E)6060<�ǹ�Z6;6;6;;;;;;;;;;B;B;BnUBBBBBBGBGININVNNNNNGNGNGNNNN<iVGNNNNNN1���V����������������tL������������������oDa�˻����������������������B�Z����q���M�����������������������a�����w;BB6aNa666-!<VQ7%%)B���Ҽ��ho>����˵��������������ҁkwI���|o����������������������������`���h��Q$-03!���E000006)w���Z6666;6;6;6;;;;�;B;BBUNBBBBBGBGBGINVNVNNGGGGTGGGNGN*�NNNNNNN%�ک����������������L����ZZZZZZZZ������������˻����������������������a�h����M�՗i�����q�����������������S�����V;B66]�]06F���ڎ3)---B���Ҽ�h7�gPu����ҝoZZZZZZo����������Ji@���@����������������������������p���]����$33J��X(0-00600B���w666;6;6;6;;;;;c;;B;B;B;BBBBBBBBINPNPNIGNGGGGGGNGNG8�5NNNNNNNک���������������ė�L!4��������hQ*Q��������ڬ����������������������u�a���i���M������MS����������������S�����%B;B6;666N����N)000-0����˼h}*7uu7e�ږSz�����Ҽ�>.JQQaa���wVD���Q�������tQDMVZSJDQp����������J���i�����ݰF�ڹ!%-000000%���i06666666;6;6;;;;BMB;B;BBBBBBBBBGPNPNIGGGGGGGGGGGGBiVBNGNGNGNV���������������˒Q.*9L���������üL<<#L������Ѭ���������������������S��Z���g�՗q�����c�S����������������S����eB;;6;606F�˖{Y0000-0-����ڼhI$%!!84��F�������oa�������lX��MJ��L����oQD4���������˸�lXa����Ҡ����t����í��.�ǃ)$)-0-000!���Z66666;6;6;6;;;;;;;;;;B;B;B;BBBBIIPIIIIGBGBGBGGGGG'�!NGNGNGN<4�������������ڠL'<N?h���������˼LNN5o�Z�����Ƭ���������������������B��M��V���J�����J�v�����������������B����%;B;;;;6%�X!)00000-0-0J�����pS2jBGN;j?��o�����z]�����������ږ�}@��D��|I��`��������������ݽh]���w���J���X�~~~�@��z(0%0-0000!���?060606666666;6;6;;;;B;B;B;BBBBIBPPPIIGBGBGBGGGGGGee<GGGGGGG'e�����������ڰL'CNN?����������Ҏ=N5.����Z���鬬���������������������M��B�i���[�����q��M�����������������B���F6;;<;76-L.0000000-0---�����wZ�����4�����tt��������������ڑJ@�uZ�|�ک��������������������h��Z��o����M~~~~D��z--!---0-0!���606066666;6;6;6;;;;;;;;;;;;B;I;IIPIIBIBBBBGBGBGB*�GGGGGGGG������������Z'CNNN?���������˖8+*.o������L|�ᬬ��������������������i���Jq��՗i����q�՗i�����������������B��F666;;7;)7)6000000-0-0--i����wl�Τ>A��t����������������˭|�J}�eک�ü�������������������hS��}������Xq~~X}��$--!-0-0-B��X0000606066666666OO;6;;;;;;B;B;IIPIIBITBBBGBGBGBG<�.GGGGGGG5����������ږ'<NGNG?��������wVJQah����������o�ì���������������������B�՗iM���M����q���V������������������B�X666067!?70000000-0-0---+����w#o�h����������ˬ����oZZh�|=d�Q��X������������������������}��S�������hd~xB��/-(-----�ǚ)00060606666666;6aNa6;;;;;;;;;;BBIBIBI;BBBBBBBBBB.�<GBGBGBGGI����������N?GNGNG?�����ݠSi�������ü��������ڸ����������������������g��oX��՗i���q���g�������������������Bs-6666%X�D7770-0-0-�-----(i��õ>��������ү�~����La���˼�|d�@�X�����˱h������������������u�B��������d~=�ǚ$-!---08��/000000000606066H6]�]66;6;6;6;;;;IBPBI;BBBBBBBBBBB8�.BGBGBGGA��������ک!GGGGGGGM����S�����������ü�������ڬ���������������������J���ZE���M���q��եq�������������������B-060%e�ˠ57700C-0-0-----(-+����7�����忝~������Dp������ü�|Xt�X��������h������������������uB���������dqJ�ǌ!!$--E��E-0-0-000060606666666;6;6;6;6;;;;BBIBB;I;B;B;B;BBB.�<BBBBBGB5��������ک9GGGGGGGL����h��������������ü������ì���������������������M���4�tg�J��q����J��������������������3660Q����!77730-0-------(((qi���d����گ�~������gp�������ü���||Z���������ݬh�����������������J��鲕�����dk��q+!XǰE-0-0-00000000006060666666666;6;6;6IBB;I;B;B;B;TBBBN�.BBBBGBGN�������ک9GGGGGGG'���t���������������ü�����ø����������������������o���7Qj]#��i����c������JV�������������!60Q����e0707030-uu--(-(-((+���V����ݥ~~�������V���ک����ô�����}���ݚ�������t�����������������t�ؕ~~�����dtJ������X!-----0-0-000000606066H6666;6;6;6;6BBBBB;;;;;;;B;B;!�<;BBBBBB!�������ҩ9GBGBGBG9��钳�����������������ü���|o����������������������S���u��L_:�V����[�����q[�M�������������0Q�����!-037333Y@NY(-(-(((i��waax����ڎ~~������|Z����Z����˼��|I�������4��������{����������������X~~���������|�Q8#!!------0-0-0000000000606060666666666;;I;B6;6;;;;B;B;9�e;BBBBBBBX������Ҡ9GBGBGBGBh��h�������������������ü��t9}����������������������S���u��՗+g���՗q����J�՗q�������������!F�����h00-0�73--��--(-(-((+�ø2@N2t��鷎~�������|�����i�����˴�|�������v�ee��������e����������������tq����������D����3((-(-(-------0-0-0000606060666666666B6B;B;B6;;;;;;;;;<�)B;B;B;B7������˚9BBBBBBBBL��h�������������������ü�|29B�����������������������S���u���o����եq���Jg�եq��������������������!0-03-333(-(-(((((((i����X���~��������|�����w������í|��������S�Sc��������t�����������������=�����������L���w!-(-(-------0-0-0000000b��60606066666;;;6;6;6;6;6;6;3�<B;B;B;B3��������!BBBBBBBB5��t�������������������æa2.GBW�����������������������B���u���o���Υq��Jg��՗q���������������o�����z--0-0--3-3(-(-(((($(E��S..��ݥ~��������������w��������|���������a�{����������h����������������k����������gi���3(((-(-(-(-------0-0-0��PG�b06066666;;;;B6;6;6;6;6;3�e;;;;;;;;X�������<;B;BBBBB9��t���������������ڸwZJ*;B;!eì����������������������B����a�����²J�Jg����[q����������������{�����B-----(3(3.E(((((((($��Vz�ڎ~��������������p�������һp��������v��{h��������t�����������������W�����������Zi���!(-(-(-(-------0-C-0]ou7*�006060606;;;666666666;6N�36;6;;;;!�������F;B;BBBBBBQ�t���������������i<%337.%<i�ڬ�����������������������B����Q�¼�ȼXBg���՗J�����������������S�����)0----(3(3(-(($($($$J�ig���~��������������l���������p���������>���oz䤕������D����������������D�����������.i��S!(((((-(-(---------\)!%!!T06060606;;;;;66666;6;6N�)6;6;;;;3�������F;;;;;B;B;F�t�������������>4]]gg{{������ì�����������������������B����a������E���՗Mq������������������J�����o----((-(...(((($($($�w*�������������t�ҕ�Z����������p��������hJ���o��~~~�����@�����������������|�����������>X��.!$((-(-().*-----0Kj;NGB�000000006<;7606666666N�<666H6;6;7������X;;;;;B;B;.�t������������hz�������������ά������������������������B����h����������[i��������������������B�����!----(-(C(.(.$($($$$$P�t������������h�φ~dX���������v������孂XJu~����~~��ؕXX�S���������������t������������JS�}J!(((($.@.$-(--y---������-00000067;7606666666N�<666;6;6;-������}3;;;;;;;;3�t������������t�������������ږI��������������������������Z���ȑ���������c����iS����������������B�����!(-((((((((.(.$($($$$�*��������������҆~~=����������h������~D�Z�~��L=g���~��~x@�D����鳤���������l�����������w�h�XB($(8@*)(-(---Y---T��ߊ-0000000777006060606N�<66666666-�������-;6;6;6;6;h�����������d�������������Io���������������������������p���¼��������T���Ja��S���������S�����]����(-()$-(((($($.$$$$$$$!�Q������������tݎ��=q����������z�ǃ���~~=�az���#z@�����~��@�zL����鳖���������i�����������X�h�X3e�J$(((((-(-(---------0-0-0777776060606N�<666666666F������);6;6;6;6;Ft����������ᜨ������������vIo�ֻ��������������������������w���¼��������iqMv�΢V���������S������Z����c-((!((((((($�$.$$$$$$$q�������������Xݤ��kX~����鸆��i���1�φ~ma�h���~@���������go�1������kt��������~X�����������h�hQ`�L�V$($((-(-(--C------0-0-0007770000000N�86060666667������$666666666<h�����������X�����������zSQ����٬�������������������������i����¼�������Q`���՚V��������JJ�������w����!(-((($($?$$$$$($!$!$!h*������������tǆ��=~~����~~~1J���8��~~Q��}o���QoLL��������D�Jz�����~=q������~�J�����������X���a�e!($((((((((-(-(---------0373030000-N�8606066666$������766666666;2`�����������p���������SQ������黬�������������������������J����ȼ�������7���՗i������iB+q�������S���ݚ$((!((($($($$$($($$$!$7h7D�����������Xڝ��Dq~~���ڎ~~XX@��|J�~~�D�Q����*���������X��L���~~��J�����ҕ~��g����������M��a�X�!$($($($((-(-(---------0-030-0000-��80000H0606$������7666666666%^�����������h��������So��������ʬ��������������������������M����μ������g����[q����iJBJi���������J����8(((J$($$$$$$$$$$$!$!$!..GNGD����������XoǗ�t=~~~���~~~8�J��Qu����8Xȁ@����.oJL��������L�L��������D����������tX�������p�|X�J�Ú!$($($((pp((((-(-(-(----3330-0-<��8000060606$������F666666666-J���������کh�������So�������o�����������������������������v������h��aQ�����c���SBJv�Bq����������B��˭(((Q3($($$$$$$:$$($!$!$E�EZ���������Xs����*q~~~���~~~D�D��a}����B�z[g����LJXJ��������.��L�������t|�����������X�����e�L�øa��Ú3$$$($Y@NT((-(-(-(----3-30-0)eک8000000000$������X-60606666-J���������ږ�������Do�������z>tݻ���������������������������J��������uw����եJ�iBP����ǒ�����������E���a$($(3w!$$$$$$!$!$!$$$!!!Z��������a�XǗ�L=��~~~�ǆ~~mZ�@��a�����J�%;w���wJgJa�������wL�S��������L������������wJ����a���e���Ú�B$($($��((((((((-(-(-(3-3)8��e)0-0-0-000$������s)60606666-����������ڃ�������Xo�������tt��٬��������������������������q��������������ե`JJv�����̒������������Q���3($($$@;!$$$$$$$$!t$$$$!$>*Q�������a������q��~~~��~~~J��D��a�����B��.X����JJw�a���������7��������L�������������*��X�ÁJ�h��Ú]�X!$$$$($($($(YY(-(-(3-3!�ږ8-0-0-0-000%������sBJ%06060-����������ڃ����μ�Q�������%F���黬��������������������������M�������������ե4P�������̒�������������a���$$$$$$$7;$!$!$!$P$!!!!!*J������a��Q�Q=����~~~�~~~J��Qw�a�����B�oXȫS���oJ..Q.DJQLDD*S�DL��������L�����������i�����X����h����X��$$($($t$(:?L6(((..!e��I$---------03������s+o���C060%�����������e���μ�Xo�������N-Q����ʬ��������������������������i�������������ե:��������̒�������������J���3$($$$$$$$.�Q.$$!$!$!$$$!!J�����X���D���JJ�����~~~~~~Q��DX�h�����:ofuȼ�}�DQ.sZ��h������.*Da��������|���������i�L���XX�����X���ÇJ{e$$$$T($G��C(($e��e!(---------%X������swo����!-N�����������w���ü�S������ک%6N����լ���������������������������g��������������+��������ǒ��������������@���$$$$$$!$!$B��3!$!!!!!!!!!����s����o��ZVz������~~~~�D��DJ�hw����.8R�ȻXJJ���X�>��Xw����w.�S.DQ������S��������Z�h����@�DX���������ˎMV48!($$$YU$V���V!((-(-(-(-(!`�������X)!wwo��w4����������ږe��Ҽ��Q�������e-6F����Ử��������������������������J��������������Ep�������ǒ���������������D��S$$$$$$$$$$$!���!!$!$!$!!$!.��������a���IQ������������D��Qa�hQ����Q����h������|Q..QQ..w���JX�JD�a������h��������h���ҖD|��Q���X������Î.SVZq�iS+$((-(-(-()`��ü����B-0$`�woo+4ZI@JJ@Ii��S���ü��a�������B60%����ڻ���������������������������q��������������[J������̣�����������������Z��$$$!$!$!$!$!3��!!!!!!!!!!���J����J���Z@������������@��a�S�����h������¼�JJZJQ..QZJJJa���h��a��������>������X�����i�S���o���a�������˭i8!$!!($.$((((((Q�����ü���!----$JwBg�P|������S4��Ҽ��so�������B60-�����ά���������������������������M������������՗Bv�����ǒ�����������������S��;$$$$$$$$$!$!$��!$!$!!!!!.a�������D��Z�@������������8��Z�X�JX����o������X|Q.D.Xn�h��h�������SX�L���������S��L���L��J�����������˖iS8Vw��������ü�3)-----)!**wo��Po�������iü��S|�������B000?���ÿ����������������������������i��������������MB�����嵒�����������������B�;$!$!$!$!$!t!$!��!!!!!!!!@c.�.�����D��MwJ������������8|�QȼXaQJJ��Q������aZ.X��=�بo7@>�Xn�X�������17����������Q��L����X�a����������eX�����������������������Ҳa3$(-(-().*o�Bwo�ڎ4I|������X��Q��������!000?����ì���������������������������q��������������[iv�����̒������������������@;$$$$$$$!$!$P$!$��!$!!!'@c\U������J��iZJ������������1a�a�ȑJ.�������������|X��������>J.�J7|����i҃�������娃��wo���L��h�����������iMa������������������˖8(((($8ZIL��iBwo���iڃ|�����}JL�������L)000?����������������������������������[������������՗qB�����ǒ�������������������$!$!$!$!$!$!$!!!J�a!!!!!;p\\NGS2Q�����Q���SD������������D=����XQ.�����Q����՞Z����������>..Q1#X��`҃��������t�����=����X�h�������������ϥvhSZw����������i8!]i���e|��V�ewwo�`��eS������Q������o.-0--;����������������������������������c��������������Ji���ݵ��������������������S$$$$$$$!$!$!:!$!$Z�*!!!!'p\UNGB.�����Q�h�S@�����������wX_��ao�X��X���������������������JQ�.BJS҃������ÑQ������a����D�|�S���������������������������i���o���\`oB��e��X�����a����o.)-0--a�����t���������������������iSS����c��������������[q�����ᒒ�������������������B!$!$!$!$!$!!!!!!�o!!!!R\UNGB;7h7�����D�h�SI�����������af�J���Ȟa.a�XXJ�����������������J..niS`�I��������.i�������Q���ZQ���X��������������������������������������i����I���ږw�e��ü�X�����L�o.)((--)o����o@���������������������V�ή`��c�������������՗J������ݒ��������������������$!$!$!$!$!$7$!$!.�*!!!!8cUNGBB6GNGq�����J�a�Va�����������a|�dk�ȥs.X��aE������������t���*--�JBXw�iJ������ҭ#X=������@��������}X�����������������������������������l����w�����ږe�˼�XXJ�����XQJQZZJJ*@JJ@@o���������������������J���XE�������������եS�������ڒ��������������������!$!$!!!!!!!!!!!!|7!!!!'c\UGBB;6E�E�����M�Z�g�����������au�DJ�a�Q.hh¼�_�������������@!�Zow���J�������XnJ~XX����=����D������XX��������������������������������l�����J���ږS�Ҽ��XQQc]�����X��������QJDo����������������������`t��K2Q8�������������եS��������ڒ�������������������J!$!$!$!$!$!$!$!!]7!!!!N\UGBB;66�����V�Z�a�a����������hn�@h��Q..�`�7��¼�����������2f�Qow���Z�����t8d��J~qX���a����|��������X]�����������������������������l������V�˖S��ô�.o��ᩁ�����h��aJ@JZ�������������������������`J��tgx�Q�������������gS���������ڒ�������������������+!!!!!!!!!!!!!!!!!!!!!2cUNGB;666�����w�Q�h�J����������hJXZQȗa����h���������������8'!Y2PNHa�Mo����a����Wq~~~��J~~X���������o��������aJa�������������������������t������|�eV��æXo�������ݬX�����X*Z������ZVJMQZJ.+v����������J�T��L���u������������cwP���������ڒ������������������i!!$!$!$!$!$!!!!!!!!cUNGBB;666����ڸaJ�h΁�����������#k�D��.�����o��������������P�>��R��BoJJ��h����@~~~~���Jq~X���������Q����������XV����������������������t�������Ii�ҭaXz������������]Q����a.D*JZo�����XJv���vJJv��YBx�J��z��պ�Q���������՗J�J����������ڒ������������������B!!!!!!!!!!!!!!!.7!!!!U\NNGB;6666������XJ�h��X����������.`��7a.�����ox��������������Q֖G#��@��+X��cJ�����=~~~~~���Dd~L���������SL��������ü�VV�����������������>����������aXz��������������ҸX!D|����Q*JXahJ`���������v``��PZt�s��u_��tKo��������[q�i����������ݵ�������������������$!$!tP!!!!!!!;o3!!2cUNGBB6666%S2������.�o���X���������Q1��L�E7����rhG����������������ng\UBN��ta��JJV�i����1~J~~~~����tXXd����to����SL���������ü�aVMSSSVgggchhh]ZS����ü��.o����������������ږ!-()t�����Q@k�����������������YMx͜��z��hDtcUB?�����՗J���P����������ݵ������������������J!!!!!!!!!!!!!!;�*!!*ccUGBB;6666!�������J�����X���������h_g�|Eǥz���3���������������u��x�ttm�Qw��+���es3DMJdd~J~~~~����t1J�����t@|����XD��������������������������]������üt����������������ک8$-()k����LL�����������������YMx����t����g�.B60(H����[q���Y�����������ڒ������������������%%$!!!!!!!!!;�w!!*ccUNGBB66666w�������a�X��h`���������=dg�|�ե����t�*E�������������G������=���7���wA;�qJ~J~~=X~~~�����DX������|L������QDa������������������ü�e��������i�����������������I)(-('k��X8Q����������������YMx������j��7��u�?($$$$aaJ����J�����������ݣ������������������J6%!!!!!!!!!!!B��7!!.cc\NGBB;66666w������ݼJ����Q�#��������Xqd1gg������֓t������������Ea�7wZ���i���w8$6$J~~J~~R1Xfx�����tDz������L|�������haQJDDJJZZZZMMMMSSZS4���������X���������������!-(-(3q~X8g���������������YMx���������t��aZ��uե!$$$$$0Fi���`�����������̒�������������������%66!!!!!!X��|!*ccUNGBBB;6666%������ݼ������P�:dX�������X~~X7g����鼗�r���������ؚ����������ٚ���x��ڠXX#1~~~X#8ZZiwwZZLQ���L=������oL��������������������������e�������ˊ���������������M$-(-$=~X8g�������������vYMx�����������j�騗Z��o�ե!$(--F�T��qx����������̒�������������������i-66-!!!!!!B����*ccUNGBBB;66666!�����弼��Q��X��Bmq=X������Xq~dau����7<7�������������������������������D~XX1@D������������xLQ��Dk������LL�����������������������e���������Q�������������!(-(-'XX1`�����������vYMx���������������j��a�h��h��ե?3io�z�qp����������ᣒ�������������������/;666-!3�����>*VccUNGGBB;666666S2>�����ü���X��P��D~~qJ8Qh���>=~dE�����lJ����������������������������a���A~~1D�����������������xLQU=�������LL�������������������ҩ����������h������������M)(-()'81X~�������vYMix������������������v���o�h��a���gi���B��JP�����������ᒒ������������������i.;;6666%Q����|3@VUUUUNGBBB;6666660z����ü�����hX��4#~~~Jx~mD=a�J=d=�����E�7����������������������������V��ݥX~R���������������������x7g�������Q@o�����������������h���������e�����������!-(-$#Dm~~~mXD8Dix�����������������������M��X��h��Z�gJ�����J��>�����������嵒�������������������/B;;666-2����X!5NNNNNNTGBBB;6666666!SS���μ��������J�im~~XX~~~~m#11XdD����g�a����wzz���������������������.����8=�������������������������xDo�������o@Q��������������p����������e����������M$-()'DgmXJ@1Zx���������������������������ؗi��g��Z��7J�������i}�p����������ڵ�������������������i9BB;66-o��oJ%6BBGGGGGGGBBB;66666666>��ü��������T��+D~~xD~~~~~=q.~d#�����՞��gJҙ�j�������������������7#����ta����������������������������i@g���Zo��LDw���������Ê����������e���������e!$#8Zwz����������������������������������M��J���Zw�B��������ig��J����������ڒ�������������������3\BBB6-|�o2-06;;BBBBBBBBB;;66666666->*iü�����������J#~~~1~~~~~mJ~~~da�������E����B�������������������8X�����a�����������������������������ޜi8j�wBD|�oDDa������������������e�����ڸeZx���������������������������������������՗X�wM���7ooB�������J�+��B����������ڒ������������������i!cGBB3|o2-66666;;;��BBBB;;666666666*������������J��x~~8~~~~~~8~~~~.��������i���B����������������ୁ=xa����t�����������������������������������ͤX+o����ZDDXw�d����������h���ÐiViz���������������������������������������������aoooo՗7>ooB�����iP��S��M����������ڒ������������������+mUG3L.-66666666b�LL�h;66666666666-.�����������d��4X~~Dt~~~~~1~~~~#�������ե[���B����������������ȥ՗X=�����g������������������������������g��ӚP��iJB@DJZotZ*�����������J��Qi��������������������������������������������������BwoB�MiT�BoB����Jv���i��M����������ǒ�����������������igU?Z3;66666666buuuub66666666666a����������X��JD~~Jf~~~~~Dm~~~Dg�������եq��B��������������������U8����娥�������������������������������鱖��ì������iJ+�����������JQx���������������������������������������������������՗`wo+i��ztBoB��iP������m�B���������ڵ������������������+RN79B;;6666666�**�6666H66666.����������s�q#~~fJ~~~~~XX~~~X��������եq�g���������������������H������l����������������������������i���o������ø�����`���������騜������������������������������������������������������awwB���J�BBoo+B��������`�J���������ݒ�����������������J!#*CGBB;6666666K!K66666666-X����������i�qx~mD~~~~~fJ~~~x#1���������ե�����������������������V������o���������������������������p���S������������d���������峭������������������������������������������������������gB�wB���r�iqXoB���������`�S��������嵒����������������q.\UNBB;;666666\N%-N\6666666%S����������g��f~t@~~~~~fJ~~~~#XdR���������������������j���������ܜ�����峗��������������������������m�ƍY����������ږ���������峭�����������������������������������������������������gJwJ�wJ��J�i`BBoB�������ڼ`�S��������̒�����������������+!X#N\NGBB;;;6666O�\BB\�b66H6662.���������U��4J~~1~~~~~fJ~~~~18~~=g������ե>��������a������������Q�����鳥������������������������ww��`o���������ک����������Z��������������������������������������������������՗MJ��J��J���B�+v�BoXi��������`�S�������̒�����������������J=qX8\UNBBB;;66666bĄ��b66666%*���������U��4J~~1~~~~~fJ~~~~11~~~f#g�����¼�������g�������������ڧ������鳥�����������������������uw��Jooooo��������������ݰ�a������������������������������������������������՗Mp����B��B��`�`���JooV��������`�J�����嵒�����������������qd~dg\NGGBB;;666666��66660%@*a.��������M��4J~~1~~~~~fJ~~~~1m~~t8q#g���������ܜ.����������������Z������鳗����������������������uw��JoooooooooX���������Җ��p����������������������������������������������՗Mv������J��BiB+�B���iXwB��������`�B����̣�������������������M��~#.cUNGBB;;;666666660!c>>��������M��iJ~~@~~~~~tJ~~~~@#D~~mD~1a.g�����ԚD1=����������������Za�������o���������������������uw��SooooooooX����������\���i��������������������������������������������՗Mv�������S��i+v�X�i����Jwwp�������`�B���ڒ�������������������J���.G\UNGBB;;666660-6#5a*?L�������M��qJ~~1t~~~~tJ~~~~@1~~XX~8m~X#a��a11~~=X���������������h����������l�������������������պS��SoooooooE��������Ú4����Z������������������������������������������՗Mv���������B��J��P�B�����iwwX�����ڵ`�B���ǒ������������������qg��XNUNGBB;;6666%%!9#**��*X������T��qJ~~#t~~��tJ~~~~@#m~Dm~@=~~~=8XXXdd~~#���������������uا���������g�������������������B���BoooooT���������`XBw���B����������������������������������������՗Mv����������JB��B��X�|������BwwT�����i��S��ڣ�������������������M���w!UGGBB;;666X%%!K.>>������X��qJ~~f~���|J~~~~@8=~1~~18q~~q.~~dXdK~q=������������՗��إ����������i�������uuuu�������M���BoooXX��������XBooBw���J��������������������������������������ΗMv����������PP�X��B�J�J�������hw��\����J��i��ǒ������������������V���7L2P5GGBB;;66H-M#X����Ãx�qJ~tf����|J~~~~1#8x8~~1q=~~~==~~dKd=qqa������������o���إt���������g���go��ýj.Qo���h���JooE�������Q@BooooXi����g������������������������������������gJv����������PP��pw��B�X����������J���BSZS�w��ڣ������������������J���L�u}!GBB;;66-M����˚`��J~fJ����uJ~~~~1RGJ~~1~8x~~qq~~d1K==d������������Z������o����������eaZ������ڧ���aQQw���+L�����Q@BooooooooB����J�������������������������������κoMY�����������PP����S���J`�T��������ک`��������J��ǒ�����������������q|��|�GBB;66%$`X���˼S��4J~JJ����uJ���~8Gq~~qXX~~~=.~~~~X=q=1�����������a������՗az���������iV������ا�����T�XL���ZDBJwwwwwww���wXi����V��ȺuuuuuuuuohhhhhhhhZZZZZZZZMJ`������������PP������e����������������کi������w��ᒒ�����������������L��|*GGGB66�B3�����\��4J~8Q����}J����#88~~t1D~1~~~qX~~~~q=~X#��������՗�����������oaz�������ږVa���Ƚ�����QDDBXwwwwwwwwwwww`BB+�����w#8JfgN1#DZ}�������������������������vP��������w�����\������������]����w��壒�����������������M��|@UUGB;0)`X����e��4m~#Q�����J����#J~~m@1~XX~~~Xq~~~~q=~q=��������a��������������uaVw�����˼�haZJ.8XmfJJJm|gZJ@#11@@DJJXftfXBBJB:mfD#*DZz���������������������������pB�����������J���r���������������tBBB��ᣒ�����������������V��|\cUNGB%S!Z%..���Қp�4S~mQ�����Q���nm~~fJDm~1~~~~#=~~~~~q=~m7�������a������������������uohZQJQZJJZo��Q~~~~~���������oQ88DXffftttffaN1#@JZ��������������������������������Pv������������p��r���������������������̒������������������J��|ccNGGB*;h7$3Qa*�����P�J21~Da����og���Q#~��XXq=~XX~~~XX~~~~~q=m.�����ΐ��������������������������������էK~~~~~�������������oZZZZZZZZZZZo�������������������������������������Y���������������ww��������������������ᣒ������������������`|�|*c\NNGG*ho-f*F����\�qD~#a����Zu���QD���Dm~8xx8~~~~=q~~~~~=K�Q�����Z���������������������������������է.~~~~~~������������������������������������������������������������Y������������������������������������ڵ��������������������i|�o2�Zuppp*J�LL�JU%���ږhXmw����X����Dz���8~~XX~8x~~~q#q~~~~~#�a���ȉ�����������������������������������է#X~~~~~����������������������������������������������������������P�����������������������������������ڵ���������������������qt�718]Zc\GNBBb>uuuu>7b-e����Jq?2?x=!�����Q����*#����8~~x8~XX~~~~X#~~~~~=������X������������������������������������ا=1X~~~~�������������������������������`J������������������������P���������������������������������ڵ�����������������������@LD8<xcUNGGB*o**}!-u4����e�+ouo#q<3�����D����Q���uJ~~~8x~1~~~~~..~~~X�������a�������������������������������������ا=X1X~~~~������������������������uQD88X|̥����������������������o������������������������������ڵ�������������������������+Lo*1tcNGGBB*7!D!B=%����p4S2hS2X=)(!�����D���}����Jf~~~XX~Dm~~~~q.~d���������������������������������������������ڧ.qX1DXx~�����������������oQD11@Jft~~a��̞����������������������o������������������������ڵ�����������������������������+7�L8ncNNGGB*YN%-NT-\!b����Tim!.�����D���Z*����#f~~~x8~mD~~~~~=.��������h����������������������������������������ڧ=qxXD18Jfu|��kQJD811@DJXmx~~~~~~~a����ܵ�������������������������������������ڵ�������������������������������������+*oDnUNGGBB*7�\BB\�>$T#%#����B>*+8=Q�����J���@Q����m~~~~8x~1~~~~~~.��������������������������������������������}��������H.=m~~xfJD@18811111@@@@@@@111111U�������ڵ�������������������������������������������������������������������������+1.anUNGBBB%J����J!<D%�����]+*59!KkCa�����Q�������Ltd~~~XX~XX~~~~=g������¼�������������������������������������Η�������ܜ181Xx~~~~~~~~~~~~ttttttfffffKj����������س����������������������������������������������������������������������+81gnUNGGBB!Soo!-U!#����`B>���>.H$!#=�����a|��z#����t8~~~x8~x8~~~_���λ�oooo��������������������������������������Υ���������UXXD1DXm~~~~~~~~~~~~~~~~~q=��������������Ⱦ�������������������������������������������������������������������+*=Qt7tcUGGBBB2I#!���˫BJu%1uJN>(8!�����Xu��Qg���L~8~~~~8~~=q~Q��������˽�����������������������������������������g����������DX~xXD11DXx~~~~~~~~~~q=j������������������ȕ���������������������������������������������������������������+88DJZZ�����LxcUNGGB;.Q-#�ݼ�a4�7�7�RU7!%!�����Q���D#����~Jm~~~Jm~q=X�����������������������������������������������������g�����������DXx~~~mXD18DJfmtfX8j����������������������¼������������������������������������������������������������Eu����������L1tcUGGBBB.\%�ݼ��=8..8#X<$%!!�����D���8X���D~fJ~~~fJ~~88����������������������������������������������������՗�������������i8Xm~~~~~tfJ87�����������������������������¯�������������������������������������������������������+Xfmqx�u|�Q*8tcUGBBB;aa�:3%#ü���*D$ITnI(%!!�����*���x~��1~fD~~~x8~~XZ������������������������������������������������������Z�������������ޜxZ11@@11iz����������������������������������ȴ���������������������������������������������������+DtcUGGBBB%2@N2J!Ckü����N7-7N�z.!%!!!$�����#�~m=~~~X@~f8~~~~1~~xa�����������������������������������������������������՗���������������������������������������������������������������ª����������������������������������������������+Jn\NGBBB;%��+g+9�����=J�p\p�U!*!!!.�����1~~Jm~~~#J~f1~~~~Dx~~D�������������������������������������������������������a������������������������������������������������������������������ȳ����������������������������������������qfn\NGGBBB%+i9!=�����J�ĥQ!!!!S?D�����@~~8#~~~mm~f~~~~XX~~D�������������������������������������������������������a������������������������������������������������������������������������ξ���������������������������������`nn\NGBBB;%+i�Pi!o����Q2O.!%!!!J����uJ~~D~~~=~~m~~~~x8~~X���������������������XX��������������������������������u������������������������������������������������������������������������������������������¼��������������`xj\NGGB;;%+i��4.C�����#!0(!.!!!Z����`X~~f~~x8~~tt~~~~1~~xa��������������������θX������������������������������պu������������������������������������������������������������������������������������������������������4SVZw{xcUGGBBB04���4�����!-(!!!%!!o����Qf~~x~~XJ~~tm~~~~Dm~~=������g���������������Ή�����������������������������պu����������������������������������������������������������������������������������������¯�������������+4SZS>F�������pGBG��Si���:.����o!(!!!!$2!|����Qt~~#~~~Dm~~tf~~~~XX~~qg������Z����������������g������������������������������u���������������������������������������������������������������������������������������ȯ������������q`�h4i�������l>e���J4�������������ڻ�����:J����=%!$!!!!$!#8-!|����Qt~~1~~~#~~~tX~~~~xD~~~d�����ե�����������������g�����������������������������u��������������������������������������������������������������������������������������ȯ������������q�����www�������������w������������������λ�������:Q����%!$!!!!!$(!D%%!�����Qf~~8~~x1~~~tD~~~~~1~~~~d������g����������������g���������������������������պu�������������������������������������������������������������������������������������Β������������J��������������������������������������û���������vZ���w-(!p!$+%!t!!�����`X�~@~~X1~~~~1~~~~~DX~~~~d������g����������������g��������������������������պu������������������������������������������������������������������������������������Β������������T���������������������������������ݻ��������������:*a!J���Q-)!!!!!$T!!�!!!!$�����}J��8~~J8~~~~~~~~~X8~~~~~=g�����o���������������j���������������������������o������������������������������������������������������������������������������������Ւ�����������q`�������������������������������ι�������������`J%*%.*!J���=!!!!!.3*=�!!!$$$������@��1~~J@~~~~m~~��ux~~~~q1Q�����g���������������g�����������˼�������������Z����������������������������������������������������������������������������������ռ������������`�����������������������������λ�������Y`SJB**%**3;;6!.S#���#!!!pP(-Q�-$$$$$������8��8~~J@~~~~X~~���X~~~~~=qXg���Z��������������ؗ�����������ô�����������՗����������������������������������������������������������������������������������ժ������������]���������������������������λ������`JDDaxnjGGBBB;;#K#2!���%!$$!!!$)u�%!%������8��Lm~J8~~~~8~����*#~~~~~q=~q=��a����������������g�������üü�������������g���������������������������������������������������������������������������������Ò�����������it��������������������������ΰ�����v@Q������hQ2GcNGGB;;6=X-a.o��!!!!$-*��*������D��|J~J1~~~~#x����LX~~~~~Xd~~dD7�����������������g�����í�ü������������g��������������������������������������������������������������������������������Ւ������������]��������������������������ΰ�����v@Z�ZZZZZaa����3*BBBB;0#DK#3-(*=�w!)!!!!!!-;$=��D������Q���8~J1~~~~8X����`#~~~~~~D~~~~1����������������ե����ռ��å����������ե�������������������������������������������������������������������������������ռ������������Jt�������������������������θ�����v+*81Qh��a3%006JDJUX#.7$�h!3!!!!!!!!!Q��Qo�����a���DqJx~~~D8�����X~~~~��J~~~8�����������������ե����ȴ������������՗�������������������������������������������������������������������������������Ò�����������Jt�������������������������θ�����v+ho>.`�tjD1JakJJJZZZZJJJJQ@D(%�h$*!!!!$$o��|Q������a���=JX~~~J�����D#~~~����Q~~@������������������ե����­�����������g�����������������������������������������������������������������������������ξ������������Jt��������������������������Þ�����+7�gPu�~xncUNGB;.%@@N.a.Qh$-!!!S2����=������J���a#~~~mg����|=�������Q~8�������������������եg���ȭ��������gg����������������������������������������������������������������������������ξ������������Je��������������������������Þ�����v}*7uu7D�tjcUNGGB;B6!.B3*1h3!$-����.S2������Q���L=#X~~~*�����*q�������Q1����������������������gg�������Ηag�������������������������������������oQJQZa���������������������������������ξ�����������iBi��������������������������Þ�����v+I$%!!8.�xnc\NGGBBB;;!%h$(*>>#����|�������X���8>*#~~~8o����o=��������Qz�����������������������oZZhhZZo������������������������������������՗Qa�������������������������������������ȯ�����������iBi�������������������������ڻ�������:jBGN;j?=�xjcUGGBBB;;6.{!%h!!0?Lw����..������X���*.**X~~X*�����*k�������ux�����������������������������������������������������������������պg��������������������������������������¯�����������JBv�������������������������λ�������vZ�����`~tccUGBGBBB;;q!%l3*��*J���Ú�������X��Z8d~~#o����h*��������i�������������������������������������������������������������������������������������������������������¯������������JD@Y������������������������å�������v+Sl�Τ>*�xnc\NGGBBB;;-!h$*>>�����].����������@#~~X*�����*o�������@����������������������������������������������������������������������������������������������������¯������������J@Q����Q@Y����������������������������v+2`�xjcUGGBBB;B60!!!w3Q�����>]������X��*##.��*g����t�������Q�����������������������������������������������������������������������������������������������ȯ�����������iJB1DQu���������Q@Yv����������������������v+>>7h7*�xnccUGBGBBB;;6q$*�!H%!������4�������h�|#*.�|�����k7������o��������������������������������������������������������������������������������������uuuuuhaaaBBBBB:8@11@JXm~~~��������������oDJ`����������������vY+?LGNG`�xjcUNGGBBB;;6%.!2a%*�!!C$Y>������X�������h�*ww7�t>*7�����Da������L�����������������������������������������������������������������������uhZD1@81#18@JJfffffttttx~~~~~~~~q=8Xx~~~~~~����������������ZD@BS`v�����vYB*��*E�E*�xtccUGGBBB;;66%!$J�H!2�����ږ��������h|��*7�7*.�����7|�����o�����������������������Șo���������������������������������������oaD811ft~~~~~~d=q~~~~~~~~~~~~~~~~~~~~~~~xX81@Jfx~~~~�����������������J@!'!>>`�xnc\NGBBB;B6;6!!!S2a�!62%#������4��������Z��X>�..~���z*������L���������������������Θ��uaQau������������������������Ⱥ�uoaD8DXmx~~~d=~~~~~~~~~==q~~~~~~~~~~~~~~~~~~~~~~~~qD##8Jffffxxxx|uuuhQD*SxcUN#*�xtccUGBGBBB;;60>*!!!$��!J%!-.�������������ږ>�����.~��~X*�����|��������������������Ή������κuoaZZZZZZZhhhhhaZZZZZZ7#8DJft~~~~~~~~~~~~=d~~~~~~~~q==q~~~~~~~~~~~~~~~~~~~~~~~~~mD#.�n\U5.`�xnc\UGGBBB;;660!*!!0$˵H#%>�����]���������F>���>��.~~~~#7�����|�������������������R@D�����������������������������՗=~~~~~~~~~~~~~~~~~Xd~~~~~~~~~q==q~~~~~~~~~~~~~~~~~~~~~~~~~~m=�x\\N!h7�~tjcUNGBBB;;6660$!<!-*aAڵ!!(RB*%*#b���˦��������ږX���>>�>#d~~X7�����o���������������՗=~~~XD������������������������������UX~~~~~~~~~~~~~~~~dX~~~~~~~~~~q==q~~~~~~~~~~~~~~~~~~~~~~~~~~q=Q�cUUGS2?2?��xnc\UGBBB;B;;60-.$3?0*w�e%V#=1�����.F���������F����>��.=~~#7�����D������������ΗD@1Xx~~~XD����������������������������ښQq~~~~~~~~~~~~~~~d#X~~~~~~~~~~q=8X~~~~~~~~~~~~~~~~~~~~~~~~~�zJ#xjUD1!Zo��»�oZJouoD�xtccUNGGBBB;;660-h-)U7#��!@D%'#1#����J���������>����..��#dDq*����*�����������g#X~~�X88X~~~XD�����������������������������j=q~~~~~~~~~~~~~~d==q~~~~~~~~~~xX1Dm~~~~~~~~~~~~~~~~~~��������zJ#@R23h���������¼���Qh�~xnccUGGBBB;;66606?2?.Ss�eQ�J'#*S���De��������>.������XK*���M��w��ZoaZDQ�gX~�����h8Dm~~XD�����������������������������j8X~~~~~~~~~~~~~dd=X~~~~~~~~~~~~mD1DXx~~~~~~~~~~~~�������������g#D�������������¼�����o*D�xtccUNGBBB;;66600%ouoZ(9#��!�gZ^�=X*-�˼QF��������>����a��=*o�|@L|ZZ��������k#`�������78JmXR����������������������������ޜDXx~~~~~~~~~~~ddd1X~~~~~~~~~~~~~xXD18DJfmt~~~~���������������Z..Qh���������������¼�������o#*�~tnccUGBGBBB;;660-!h7Z7!a*s�F%%�*7�7*�**'4˼Q@V������˳.���D.��X*##*a7���������������k*`������L1.g������������������������������i=q~~~~~~~~~~dK~X1X~~~~~~~~~~~~~~~~tfJD@1111118@DDD@@@@@DQa�������Ȼ�uuuuuuu��¼����������D|�xtccUNGGBBB;;66-*8Jfn|z|gJ@S7�*S#ǖ!7Y1YD%��Q@�@�����üQ���D���a*1L��������������d*L������L7�������������������������������j=m~~~~~~~~~dK~~X1Dm~~~~~~~~~~~~~~~~~~~~�������������������»�hQQao�����g7.a�����������z=|�~tccUUGGBBB;B6-*X~~~���������Q2+�Z2s�*$)P#!GDQ�D)$@�DB��ü��X��J���J#da*L������������~d=o����t*E�������������������������������xDX~~~~~~~~d=~~~mD1Dm~~~~~~~~~~~~~~~~�������������������aJh������������ȉXX����������~q.��~xtccUGGBBBBB-#8%!#D_��������7Hϭ#�*p3!$7p!!%C#1�D--J�JB�����J��Q���amX**h��������~~~q.*o����7g��������������������������������DDq~~~~~~q=~~~~~mD1DXx~~~~~~~~~~����������������hQJQo����������������¼�Xt��������~~~X#���xtcc\UGBGB3%#6-600*Q������.t�M#2�pNBNp�!$?�.%--!J�Z;����||�Qa���J�7*Q�����~~~~~~XD���7g��������������������������������j=q~~~~~q=~~~~~~~xXD1DXm~~~~~~�����������ZZJLh��������������������¼����Q7�������~~~~~X1JXnjccUNG<'!!3666000L�����#��*G##�����@%>�*9-!!J�ZQ���|Z�8a���*SD��8Jft~~~~~~q=D��.g��������������������������������j=q~~~~~=X~~~~~~~~~xXD111118@@@88@@@@Qa������������������������¼�������Qg����~~~~~~~~xX8%!*%%*7B6;6000-L���g��*a%#2$>u>!N%%)1t@J7)Z�����|Z�8Z���D2=��D#18@DJXa8#7��.���������������������������������jX~~~~~X#X~~~~~~~~~~~~~~~~~��������������}aJQQZahaZZZag����¼�����������7#Xx~~~~~~~~~~~~xN1%.3BB;B;;66000-*|��#���+%!<*!%7@*ZU7-Q��L��zJ�*h���Z*���#18@DQQ�d1@#7��������������������������������Dd~~~~q.#X~~~~~~~~~~~~~~������������}Jh������������ȳ�QJa�������������D8XfftttffXD'15BGBBBBB;;666000)k�D���7!!-5%!!)'@NWB-J�����D~u���|���*.~##@1817���������������������������������=~~~~~.#Dm~~~~~~~~~~����������wLZ�����������������¼�X.a���������t7@8@8J@@\\NNGBGBBB;;6660000!dX���Hh>*!;%%0173!f��g�xDXu�������o=X*`�uDg��������������������������������Ud~~~~X#Dft~~~~~���������QJ��������������������¼���QJ|������kE���xxncc\NNGBBBBB;;66606000Z���t?2?*%!3')%.];8!x�o!!Q�m18|��������*d#*k��`*E���������������������������������X~~~~q=1118@@888@.���������������������¼������**Q�����X.���xtjcc\NNGGBB;B;;6;606000-#����ouo!$7%*fZ-##!#~~ZJ~f1u��������**a#XL���o*��������������������������������Q~~~~~q=.|���������Ηo7*!%%!!JZh�������.#g��~D��xtjcccUNGGGBBB;;6;6060000)���hS2B!CP-!1!8~~@J~f#f~���#����D##*|���|*���������������������������������aq~~~~~qJ8*X���������Η7t\NGGBB7;*7Z����.q~q7ttjcccUNGGGBBB;;6;60600-00���B!!-5!CP-!##J~~1J~J*X~~��1*����Z*8L����QJ���������������������������������jd~~~~~~~~tfQQQg���������²a=cUGNBBB;;;;)*o��.>�Dd~=gjcc\UNGGGBBB;B6;66600-0--����M+*a!;9B-!8$!f~~#9-J~D*D~~~~@*a�����>*8*�����.���������������������������������d~~~~~~~~������������.R\NGGGBBB;;;B#t~.>���_dq2cc\UNGGGBBB;;6;66600-0--!t���^`*7'-%3B-!1!$x~x*GD(J~8*a1~~~~D�����*8Q����>g��������������������������������=~~~~~~~�����������}.mUNGGBBB;;;BB.=qL���xtUd8U\UGGGGBBB;B6;6660000---!H���HX+(7%9;-!8!!#~~f*N<(f~#x~~~J�����*8>����|E���������������������������������a~~~~~~���������S1\UGGBBBBB;;;BG.XL���xtnccG#<UGGGGBBB;B6;6660000--(-+���^`>*7%---1!!$D~~J($!tXX~~~mo����D*a1>�����.���������������������������������UXx~~~������oD+x��tD\GGBGBBB;;;BGG9=7���xtccccU?GGGGBBB;B;;6660000---(-����X`S*(%--$'#!$$$$X~~8~J8~~~~L����Z*>>*7h7@>�����DD���������������������������������8JfqtmJ=i������JNUGGGBBB;;;;;BGG?*k�#Zxttccc\UUN!BGGBBB;B;;6660000---((!��ڭ�B2-%!!!1!!$(-x~x!8~J#x~~~8=�����?La*GNGoo##>����LXXD�������������������������������*+o��������>cUGGBBB;;6;;BGGGGC@Z���Q#jjccc\UUNG!*GBBB;B;;6660000---((-t���4J�$##!!$$-%62~~XQ�J1`���J*�����*��*E�EJ�LL�J@>����*.qXD�������������������������������7+ooB+>���tUGBBB;B;;;;;BGGGGN\\gnj@\c\UUNGGG*m*BB;B;;6660000---(((-H���W-!��